5|4|3|2|1|3|4|0|6|6|-1|6|6|6|6|6|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|6|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|12|12|12|12|12|12|12|12|11|10|9|8|7|9|10|13|&False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_True_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_;B>10<False}False}False}False}False}False(3580(3600(300^