5|4|3|2|1|3|4|0|6|6|-1|6|6|6|6|6|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|6|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|-1|12|12|12|12|12|12|12|12|11|10|9|8|7|9|10|13|&False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_True_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_False_;B>10<False}False}False}False}False}False(3580(3595(295^iVBORw0KGgoAAAANSUhEUgAAApgAAAKFCAYAAABoeZmMAAAAAXNSR0IArs4c6QAAAARnQU1BAACxjwv8YQUAAAAJcEhZcwAADsMAAA7DAcdvqGQAAPp7SURBVHhe7N0HuBNV+gZw14Ji17WLXbGi0jsKiKKCKFLEggp2KYogil3EihWw7NrLqruuXSx/dy2rrnXtDRV7w4b0es8/3yRzc3Lum8mXKcnc6zvP8yPJZCYz855D8t1kyjIzZ840rgULFpglS5YQERH94clnYpwWLlyYeosWLaoXFi9eTDFBfT+KOgWmdH40IRER0R+ZWyiGhQq6tEHFXBqhQonCQX0+ijoFJlooERHRHx0qFsNABV3aoGIujVA7UTioSIwilgLznHPOMSuttJJZY401zJprrulp376910nR9JX0448/mldeecUzY8YMOA0REVEpc+fOhQVjudxiLo1QMZdGqJ0oHFQkRhFYYD7xxBMee5zrf//7n2nbtq3ZZ599zPDhwz0TJkwwgwcPNgMHDqwdF0ReA712HIYNG2b69u1r+vTpY0aPHg2nISIiKmXWrFmwYCwXKujSBhVzaYTaicJBRWIUdQpMu+H8AlMGe7xvzpw5ZtKkSV7xdvPNN9fq0qWLmThxojnjjDNKkmnlNeS10DLK9eCDD5rZs2fXPu7evbv57rvvzJdffml69uxZO16meeihh2ofExERBfn1119hwVguVNClDdr+NEKFEoWDisQoAgtM4Q/uePHGG2+YtdZay1x33XUF49977z3TsmVL06JFCxV5DXkt+zXCGDdunOnatav3jerbb79tHn/8cbP99tvXPi/3n3rqKfPuu++adu3amd13390rcu3XICIiQmQ3K1QwlgsVdGmDtj+NUKFE4aAiMYqSBWaQW2+91ey2227mP//5TyTyGvJaaBlajz32mOncubP3n1d+cpcCcsSIEd59f5rXX3/dnHDCCaZNmzZeQSvTyjwyr/1aREREru+//76gUAwLFXRpg7Y/jVChROGgIjGKOgWm3cH8n8jtcbbVVlvN7LnnnrGQ10LL0JKdrzt27OgdzIOeR15++WVvHpkXPV+eh8xRyyxjljnqIfDcQvPBxHZmmWXamYkf1H0uVh9MNO2SXM5DR2W2I7OdGe0mflB6vK3ENF5G7SaaD5zxtc/l5l1mmaPMQyXGF/PQUcuYox6yx0m7OXnJenrtCJ7zRcnZm9df54wi25yoFPeTom2q6WM5dfpSGfNm5f4/W/L9JqBflFRiXvaNuuMtUfpGHO8hX3/9NSwYy4VeO21QMZdGqFCicFCRGIWqwJTBHu9r1qwZHB9GHK8lP33Lz+P2OPnP/P7773vc/9itW7f2fs63x4WX/eCQb07rvjH7H1ZJvGlH+bArlyzLfwO2l1tsvK3UNDIuk1GRD9S6hWHw+KLkg8j+IyD3gW5/KMkHTvZxsW1xaafLAB/eDx0V/KEWjzLWMTJZVth+UqRNvdxKz5slz9t9SbfcQs50ZS0/SMC87Bsl843SN+J4D/niiy8KCsWw0GunDSrm0ggVShQOKhKjCCwwhT+440XaCsxHH33UnHTSSbWPP/74Y+90SXIUuZD7Ms5//thjjzVPP/107eNosm9sRx3lFyfWc15Rc1TRN75oir+hxs4pzmoLsWLjc489JaaRx0dNzHxQFC0wi31olLnt8mFkLaN2ubXr9oGZWPtHgjZb7XTy2mUWxLGpJ/0kA7Up6i9oXv+5gr6kXG4hNy/7cZQsi83LvpF034jjPeTTTz+FBWO50GunDSrm0ggVShQOKhKjqFNgov8Mxey0005wfBhhX0uOEJf9KuXgHjmI58033/TGz58/3/s28b///W/ttHJfikx5Th7LT+QyT7du3cyJJ57ovZY/bfkeMkPlTfp9uR1qHqod/362YPHGy21u/PvyV7f/s8wyZuhD/rT+/ZyHhnrfxLxfZx5Zhrxm/jWWGfpQZh57Obn7D+Xnk9d+P/MG7M/TbmL2m92662RvQ5bMVzC9rFtmmcXG2+tedBq5L8uV+3Lrb6u93blc6q5zsfFB/Paw79tt5t4vzC+/DD9nuc2vQ8E21Y7PvZ43rm6utoeGgteK3I5oHf31j+P1c+NzovSTYm3qzlv7uGDeDFk3eU251fS9oux8MgrmKXwOt5ko3Jbs/2s399w87Bu4jQraN0rfwPMWH4999NFHcHy5UEGXNqiYSyNUKFE4qEiMIrDA9H8it8fZkiow/f/sNnta20svvWQOOOCAOsWh/PQt31ra44SMk+fscd9++633GvJa/rhy1iEr/6YsHwTZD5OM2g86903bmcZ/ruCDzH4te/7sdNk3Q2c8WE7tm6y8duZx7Zuo99j/ECj2+rnHGVE+HIpO473B55Zbm1Xu+doPB5u7vaXG11WQaW4ZDw3NzVu7Xrnn6+SH8nKX7TzOzOdtu719GZJJtm+h9XZfP2o7Bq1jHK+fe5wRpZ/UPuexllWwDtmiwHutgnlxXyre93KPoVwmtfxl+8/ZWaLx1jrCabLP132fyD5m38iO926tXPKsZRWsQ7G+YXO3t9T4PH9Xq6hQQZc2qJhLI1QoUTioSIxCVWDKYI/3FSsw77//fnPDDTfUGS/j5Dl3vHBfK//GHlzYSVG43377eee5tMcXKzClkHQLTJlXXsMuMIV2HbKsNyfrwwIWiPJ8wQeWO531hu2/QXrz5NfH431Ium+K9uOg55zHRV/fnzbEh4P/OEM1r/MhW4xkVfBaJcbX4a+ftZ7+ehSupzZbZ7piWYJ2rzOvrFPtfEVeP+hxPe8nLrtNZf7sMtuZoZk/CApeK/d87TirL4VZbp0MvO0ukhdqM9jWIjtvO7f4hNMrluNOE/S4aNsFvUYcr+9PW72+4Qr7HvLOO+/A8eVCBV3aoGIujVChROGgIjGKkj+R+4M7Xuy44451xslO0E2bNjWdOnUyf//738306dM99957rzdOnvvqq6/qzIdeS94w3HEuOW3EqFGjvCPRt9tuu4KfyOXncM1P5DKvvAY6BYVmHbLsN97cNynys1JtweS+ERcrMPNvwgVvuiU+sPAHQNBzzuOir29x3vRr16/Y+NxjD5xmYmb5zgeSKFFk2llpxtch25pZxkOZdaidXsYNnZj/BsybVputM526rZxxBfNZ38bVmS/gsXrZ9uM4Xt8SpZ849G0t61ikL4VYbt0M7G8ci+VhtVlgO2SKmMx09jrVXZ4zjn2jjijvA2HnldPeofHlQgVd2qBiLo1QoUThoCIxikj7YKKiUM4vKVf2ueKKK8zWW29dQMbJc2+99Vad+dBrleuRRx4xI0eOrH0s+8vIG7l8aynfZsp9ex+aY445xjvIx38cjfPGK2+Y8kFS+ybpvmlbb2TuG7M8bjfUDM3Iv1ln56n7pusst85yij2Hpg3+671wPa15i42XDPxisdg03uMcb7tz09vzutMUmxeNh7LFQv5bIJHd/uCfQu3Hxe77j3GW8sFZdBl18gp6/WKPiy271DxRX99SrK2LjS+3re3pg+YtyLJE36vDma5gXYqse8E02T4W1A5SzNjPs29UsG+geYuNt7z22mtwfLlQQZc2qJhLI1QoUTioSIyiToEp3+75/J/I7XE2KQrdcR988IF3qqAXXngBkuc+/PDDOvOh1yqXFLdSRNrj5s2b552+SMh9+zk5TZEUu/a48B703hQve89//J65LFMgPljs+fcuy7yZ+d+02PMJmTczfuiD1riMgnnyzz+Y+aDKP7aX465TicdFXr/Ag5k37dzzQx8sMV7GtbvMvFdqXp8s35++YF5Zz9w6FcxbbHxp712W+TC31y3Dy7Fgm4PyKnyusA0y44KytHIQ7S57L/dcrt1lvPcHBl5Wycf1up/IsvKvjdva+n9VMK/F7kui2PoUVbgehf9H7TyKtVnd18guF8xbZD0F+4bdvrKs/GuX1zc08zrrA9i/iEWBCrq0QcVcGqFCicJBRWIUdQpMKcJ89j6Y9njfDjvsAMePGTPG+zm8Q4cOHjmZuTyWq+bIc2ieYq+l9dtvv3nFq/yFiZ5HXn31VW8emRc9T0RE5JMrz6GCsVyooEsbVMylESqUKBxUJEYRWGAKf3DHi6hFoS3qa8nBQ3Jt8Tlz5ngH68i3k8OGDSsoOOUqP8cdd5xp1aqVN41MK/PIvPZrERERuZ599llYMJYLFXRpg4q5NEKFEoWDisQo6hSYctlELTmoBo0PI47XOu2002q/OZWfvuXE63IQj/+8LOPxxx/3npNpZFqZx34NIiIi5F//+hcsGMuFCrq0QcVcGqFCicJBRWIUDarAFHKgj70d8g2lXD9WjmTv0aNH7fjff//dPPzww7WPiYiIgjz55JOwYCwXKujSBhVzaYQKJQoHFYlR1Ckw5WdjLSkK0fgw4nwtm/wkLkeu9+7d25x88slwGiIiolIee+wxWDCWCxV0aYOKuTRChRKFg4rEKOoUmLNnz1ZbbrnlzMorrxwLeS20jKjkJOrPP/+8R77JRNMQERGVIr96oYKxXKigSxtUzKURKpQoHFQkRhGpwCQiIvqjKHYlunKhgi5tUDGXRqhQonBQkRhFnQJTzJo1i4iIiCz/+Mc/YMFYLlTQpQ0q5tIIFUoUDioSo4AFppCDYIiIiOh3r8BExWIYqKBLG1TMpREqlCgcVCRGUbTAdP9yIyIi+qNChWJYqKBLG1TMpREqlCgcVCRGsUzznXc0RERERERxYYFJRERERLFigUlEREREsWKBSURERESxSrTA/P3jxyiCxy4eSiGhPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgPWiwPz1g0fMAzeND/TJi3fBeYVmft9Xr/0dvob44a374Ty2oPnLhRowTv88/3A4vpjLT+ht/n7OYfC5tEF5kh7KNC0evWiIBz2XBijP1Jj2eBZ6LiVQpqSD8ozT92/9E44v5v/uuTzWz8SkoUzDeOTCIWb80J6B7jrzYDiv0MzvC/pMvn/84XAeW5yf6W4NWC8KzO/evM/86U9/Mssss0xRd1wzDs4r5D9Fqfl9T959GXwN8db/3QjnsT11z0Q4bxioAePUdJN1zbG925mHLzwSPm+7btSBZo1VVjLH9GoHn08blGe1/fbho+aWK8eaA/bubPbavbU566TBqX3zRZlW29iDu5rtNl3PrLD8ch65L+PQtNWE8kyD2Z8/Z2qWLPTIfTRNGqBMq03+oJG+1nnnLUzr7TYxg/dsmco/tlGecWq5c1NzyRnHml8+eBg+b3vlsevMOmuvYS4adwx8Po1QpmHcd/7gTM2BawTfuEO7w3mFfPlTan7fZcf3gq8hbhzTH85jmxgwf7ncGpAFpiNqgSl/saF5w0ANGKetNvqzt87yQT155AFwGnHb6QeZ9ddezZt2wz+vbh6aULogrTaUZzVJcTmgd9eCviK22HRD8+Hzt8N5qgllGhfpT+cP2ctcePTe6g/p3h12qJOdb7+OO8J5XLIsWaYsW9YBTRMHlGcazPvuTeMPch9NkwYo02qS4rJr863q9Dt5L7x93CA4T7WgPOO08w7ZHNo03868+NBkOI348LnbzGZN1vemlfe4n99/CE6XNijTMOpTgSm/TKJ5w3BrQBaYjj9SgbnzVhvWrrd8I3RQt13NA+OPKJjm7+ceZrbMFaK+0w/pVjBNGqE8q+nOyWcWZGgbuF9XOE81oUyjuiPzYdx2h00L3jgbZfpdn0yB+MAFhf3OduZhexTkhcg0aF4hry3LkGX508v7gayLrBOaJwqUZxqwwAwnqP91bb41nKdaUJ5x6tx259ptX7HRCmbMCQeZH95+oGCar1//u2m2/ZYFOd1+zekF06QVyjQMFphZ9abAXHbZ+lFgPn1v/SkwO+60eZ3133yDtWo7nHxT2WrbJnWm2X6z9TN/1ePXTAuUZzWdMfLQOjn6dtpuCzhPNaFMo7jn7EPNBrlvwZHW225SdL/KFk3r9kGXTIPmlddEfdgn6yTrhuYNC+VZDXO+fMEs+v0bs2jWd54l83/LlZfGu++Pl2lkWvQa1YAyraZDe7SAfUdsseHacJ5qQXnGab+9OtbJYMemm9d+sfLTew+ZHl1a1ZmmbfPtzcyPHq3zemmDMg0jW2AG1xwsMCNCDRiGFIilCsx9urU1w4f0hY4bvB+cB+nXazf4GmJwvz3hPLb6VGDu0XIbuA3LL7esObBLM7N32+3g89Lx49xvIwkoz2qS/ZBQlqJDq/j+r8QFZRpF0E/cvlMH7Q7nXX+tVeH0NpkGzSuviaa3ybqhecNCeVbDkvkzc+Vk6UGmRa9RDSjTapL9zlG/ETtusQGcp1pQnnE6pC/+NneF5Zc3I4860Bx50N7weSm24jw+ISko0zCyBWJwzSK/oPTt3AyS3X7QPMhuu2wFX0Ps2bopnMfGAlNRYKZFfSow9++0E9wGjU7NtoCvmRYoz2r69KW7zIbrrV0nR+nXd005E85TTSjTKNZebeU62+7qsNPmcN6tNi7cRQORadC88ppoetvaq68M5w0L5VkNC37+OFM61mQryKChpsabFr1GNaBMq0mO9pU+4vYbKSCCds2oBpRnnE48Yv86OWj12asTfM00QZmGoSkw0yKpArNLp/YsMOP2r79fAbchDNSAcZIjIdE2aMi3nNIxLzl2X2+fTPmmSG4vzTyWN2Q5zQJaZqWgPKvtf0/91fu20n/j2WiDdcxtV6dz3ySUqUt+Brp+1IHmzjOKn27Dp/n/u+Pm68N5D96jOZzedsgeLeC8O2yWPdAgiKwbmtcm2yjbKtuMnrehPKtm2uNm1rQnPPO+fztXURrvvj8+bactQplW219H9/e+rfR/tlxnjVVSuS86yjNOcuYL9/+PlnzLKT+lT73zEm+fzJsuP9W7ffyuS73TDMrpBNEyKwllGkZ9KjCvOHE/uA1h2PXfPnv1qD8F5nKZggaFkzb1qcA8br/MXxhgGzSWW24507JlC3PQQQeZkSNHmlNPPdWMGjXKDB061HTr1tXsusPW3k+P8lN6NfbXRHmmgeyHdPk5J3inKfrxncKd49MEZeq7ZexAb/9d+SPD7w+yL9q5R+4JpxcbrbN6Qf9BurfAB0z847zBZuN11oDziCbrrmHuy0yD5pXXRPPYZN3QvEK2SbbNn1a2WbZdMkDTC5RnGvAgn2jkfeyEPh280xQFHZRWTSjPOF121nEF/3fKkf3MaAk/M7p372bat97VHHtYb++n9Grtr4kyDUMKzPrypVhSBWbXLh3rV4EpfxFIJ02jZZfNftj++x9Xwm0IAzVgnPrtlj8isFwTJ040NTXFf35bsGCBeeaZZ8zw4cNM6x23MhOO2ruihSbKs9rkL/RxIw7N9JdsX+nWqUXgBQKqCWUqZKfxNVdtXKc/CPl2Z+SBneF8h+9Vd8d/18XH7APnFXecMci0BAf7yDh5Ds0j5DXdeVxH9GwF55VtKbajvWQgWaD5UJ5pwAIzPPlFRg728YuGFttsHHii7GpBecbppKP71fm/oKX/zBhuunVubR66ZULFC02UaRh+gVkfapYrEyowRb0pMBs3Xsm8+uqrZt68ean09ddfm4033rjeFJjyk99qK69Y501AS94Epk+fbl588UVzzz33mOuvv97ceOONZurUqebjjz82S5Ysyb1tGPPDDz+YsWNPNXu33zH2I3aLQXlW03vP3FJwig/fBuuubf7xl3PhPNWEMhXNMx+s7jbYGq2wHCz45IwEu2y1EZxHyEFl7jxIux02q51H7qNpXH0zr20vyybrhM7rKqcvkm1B8/gkC3c+gfJMAxaY4ci31fYp3XyyX3HQt/bVgPKMy7QX7zRrr1n8TBCllP+ZMdYM7r+3+eLVe+D6JAFlGoYUmCuttGK9qFn+8AWmXDXggH27eaGkdZC/zA47uL/3nxBtQxioAeMgV+5B3waVS/4KQuPlL6PNNtvMnHjiiebtt/P7fb3xxhume+d2ZspJfeF6xQnlWQ3yF/h1F48ya6y+CsxKyF+5QwbtY7554x/wNaoBZSqFo+bUGbLrBZr/wQuO8L4FWts5YOKwPVvC6RH7iPJiR44j7qlmZB1knKwTml6z+4hkgfY/RXlW25yv/msWz5mR+59ovPsyDk1bbW6e1SK/uIzq38Ws0rgRbH8hfWCfttt5u3Gg16g0lGcc5DN4j87h99n3hfnM2Ldnd/PSI1PgesUNZRqGfMZ2a7tz6muW/n32Ue1Dr+XWgPWiwBRyfq1bplxkhgwZYo488sjUueLis830l++G6x4WasCo5E1Tc8qYuMgbysCBA72/XGWYPXu2GTSwX+KnOUJ5VppczUL2tUS5IJtuvL558OYL4GtVGspU/tJF6+2SbwzR/D7pg40brVA7/b7tt4fTueQnSXs5QvszpSzDn0eWXWp3jaBvPW3or3+UZ9VMe8I712WxQZ6TaeC8VeLmWQ1ypSfZ1xK1OSJ/7FwwtCd8rUpCeUYlfyQfc2hvuN1JQJ8Zhx06qCKnOUKZhiW/jFw0+uhMzYJrhmo7e9Rx5u6zDoHrHpZbA9abAtN31XnDvCsIoI5ZDfLt0wmH90nkUlioAaOS/c3QdiRtzTXXNH/729+8NwzZ12bI4YeZq4f3gesYB5RnpchlISdNGBn4rWUxst/O4QN6Vv0a5ShT+dBF6+zSXK9erhzlT7/KSo28n5TQdLazB/coWI6QcWham7y2LMOfR5aNprMd3attwXKKQZecRHlWxbTHzeK5P3v/52SQnyBff/11j/1zpEyTpiPJ3TwrSU7ML/veBn1rWYx8FvRss21Vr1GO8ozq3FOOgNubNPcz45ijhpjn7r8armNcUKZRDTugY8H7XbXJt+59Ou2YyCWf3Rqw3hWYQk5rsP46a8HwKmmlFRuZay86Ga5jHFADRnHKgN28N0G0LZUgP4Ocf/753lfzCxcuNIcM6GtuPa340bhRoDwrQb617N6p+JU/tJpstG5Vv81EmQo5VQtaX58cZa1pU/en9pP64YODbAO77lIwj5BxaFqbvLY9jywbTWeT/e7so+SRYifZRnlWw8KZX3ofzjK89tprpmnT/EmXt9tuO2+cP8i06DWqAWVaCfLHguaqUaWsu2b1vs1EeUZxw6WneH/0ou2sBPczY8jhh5j3n7kVrmscUKZxkNP3rbUaPjiykuRyuSf37wLXMQ5uDVgvC0whnaz5Tvkr0UjhtNJKKyXKP+pKyEmz4zypOoIaMCx587S/xbFVuug855xzvA+1X3/91ezfo1Mif0mhPJMm53SLshO8S97Y5dvxGe8+CJeXJJSpuPbkvoHf7mi+vZT2dufbbtP14LS2Xbeue5CQjEPT2uS13fk0fS7oW0zJQLJA86E8K23Oly95/8dk+PDDD71vg9xtkHFycIU/yDzotSoNZZo0OadllIMeXfKeKt8SFdvHNykoz7Dkj+XVV8O/wlTzM2PwQfsn8ouhQJnGRf7w3qbJOrXbVOmaRfY7j/Ok6ohbA9bbAlP88Nb9ZkDvrl545557bsERUkm4//77vWW13nU78+Hzt8N1ihNqwLDk/G1+R7PJvhjyk9lf//pX+HwSpNPffvvt3hvGf//7XzNk39JFSblQnkmRNzu5HGlSb7otmjX1jkJHy04KytQnJxyXo6/dbyHlr+O/Fjl1j+3+8YcXzOcLOvhLfrpEfyDJuGLXMBfymu48QtYBTW+TbZFtsueTbZZtlwzQPALlWWn+AT1Lly417dsXP2BJnpNpZJB50GtVGso0KfKHhlyWz+3LcWnaZN3Ac6bGDeUZlpyvF21TGj4zzhszBK5zVCjTOMn7TtfmW3nbVMmaRf7Ivn1c8dO5xcWtAet1gSlkB+QtNt3QPProo17nS3L48ssvzfLLL2++fO1euC5xQw0YFroayn777Vf74XLyySfXeT5Jq6++uvnkk0+8ZZ865hRzXcAHdhgozyTIkd9dO5a+0kxUskvIs/+8Cq5DElCmLjmq3P2WT67GE1TwCdlHzZ7HF3RNcOkfaB4R1HeKHdBWaj852QbZFnse2dagc276UJ7hTc3uH+mD0xSa9elT3uUfZXjyyScLtgGRabwhM8+sT56Er1lrWvnrUy6UaRLkyO9Sp92Kg/w0etWw5PY3t6E8wzptWN2D6tLymXH6aaeaVx67Dq53FCjTuMkBhhv+efUK1izLmXvPqczpAd0asN4XmKLplk3MRhttVHt0VFJ22mkn71sqOS8nWo+4oQYMa4Cz/9oqq6xiPvvsM68TysltV1ih8gdOde3a1Xuzkp899u3S0vuPh9Y9DJRn3L79332mTfPt4LYF+c9//uNlL2/W6Pli5OeqZ+6L7zyrQVCmiBRc7noO3bcNnNaHjgYXqzZe0TwwHv+k6O5HaSu2/6a8lrwmmqfU0eeyDe48muJSoDzLMfvz58yCXz4xS+b9amqWLvb+j/pDzZKFZsn838zCX6ebud+8liny6h4BPufLF3NTGzNmzJg62+GSK6r4g8xrv9asz5428354xyz6/VuzdOFsWYHclNmhZsmCzHr+Yhb8PM3M+eL5gnnDQpnGTa78hHadKCXs/135pv3KYfGdb7AYlGdYo44dULgNKfvMOGzAvrGfiB1lmoQm665ZwZplGdVBlHFwa8AGU2CizpiE+lpgHtB5p4LtOO+887w3CjnZapMmlcvP9cADD3jrccklF5tLj4vv1EUozzjJkeL7dm8Ht6mUL774wtvmgw/GhVYQ+SZT9o1C6xQnlGkxcl1mex3lZ+Wgn5Dlpxp7epsciIbm2btt8UJenkPzyGuh6UXQz0Wy7u5P47KNaFoE5akhhaX/07Z2qFm6yCz87Qsze/ozta8z95tXc88ac8IJ+GdOm0zjDzKv9xpfv5xZlx+9bzXLGaTYlHn9dQkDZRon+XbaPmF/OaL835VvMtFZB+KE8gxr2JEHFKx/+j4zLjFP/O1SuO5hoUyTIAUm2rYksMCMiAVmafZ5ADfccEPz+++/m/fee89ss03+QKlq2HHHHc3ixYvNzJkzTY+2uqu5aKA843T1+cPh9mhE+ZAScsLjpC+hhjItpv2OdT+sZd8zOdkwmv7mUwu/GbEVOzJ7y43+DKcX8hyaJ+iId1kHNI+ss6y7O71sI5oeQXmWIt8Sut8OTps2zdx2221m/Pjx5vTTTzcTJkwwd9xxh3ciav9nytohUwgumvm1mfXZv8ycL17IjTRm9OjRdbbFJdP4w/zMekiR6A5z5swxzz77rPnLX/7i7Tsm63PxxRd7V2Txz1doD4t+/6b0z+1FoEzjNLxvR5iDRtT/u3KBizh/qXGhPMM66uB9a9c7rZ8ZA/r0gOseFso0CSwwY4AaMAksMEvrvPMWtdsgHw7ys1jjxtU/bYJ4+OGHvTftESOGB37zVQ6UZ1zkp/F11l4DbgsiP+scf/zxtX75JfsBfvPNN9eOk58zyjlIKOnLS6JMiyl2nfHBRa7Qc8Mpxa9nLG+Gbh+QHeOXs46GdMlz7kE78hpBB27IOtjT+2Sd0fSyjWh6BOUZZP6MD73+IIOcjkWKtubNg/frXW+99czRRx/tHfAg8/iD/KQuP1f7g+ZADJkGDXJamLvvvtv07NnTOyIVzevbddddvUv/yfkK/UF+UpeCF21zEJRpXOSn8TVWCd4WWxL/d5O8vCTKM6wD9s7vlpLWz4yRI0eYV6deD9c/DJRpElhgxgA1YBJYYAZ75MIhZl3rZ0w5UMnepmqTN3EZ5K/jvrvtDLehXCjPuFx21nFwO4q55ZZbvO0LGuSDyz6lRClyXXO0bnFBmRYz4ai94TrKeSQnjzygzvRyeh80vW//TjsVTC/nkEPT2WQaex55DTSdD51iSNa12LkvZRvd6YtBeRYz99vXM62fLRDlqM++fYOzQeRIcPl2EQ3vvPMOnMf27rvv5qbODvLt6E033eRdug9NH2SHHXbwrr/sD0sXzS27yESZxkVzCVBbEv935brmaN3igPIM49cPHjEbb5j/Jj/NnxnDh/SF2xAGyjQJLDBjgBowCSwwg8m5r4K+zak2uTSYfz6+3j17xHJeTJRnXDq2Di5eXLKP2z/+8Y9ac+fO9bb15Zdfrh0nH2TlfAuyfCazT168C65fHFCmxcgR2cX61xYbrl2nPa8Zvj+c1ifnI3zAOn/g0H3qHnDjkmn86WXeUuc0lHXwpxeyjrKuaFrZtnKuzoLyRGZ9+n9GDtqRQb4t7N69O1y+1qBBg8yPP/7ovZ4/SLEYtL+cPGf/3C4/d3fq1AlOqyXfct111125VzTeQUnlHHGOMo3LTiUuFOBK4v+ufOOuvcRpuVCeYfzfPZeXtU2VZn9mHLh/b+9S0mg7yoUyTQILzBigBkwCC8xg3VtsDbclTc466yzvzeKaa64p69uiYlCecZBzXq7cWP8TGxJ1Py7fvdefA9cxDijTIBuvU3yXgYHddi2YVv7gQdPZxhy0e+30nZrld+8oRqbxp5d50TQ294TDso5oOiHbZk9bCsoTkSPB/WHs2LFw2eXaYIMN6nybeeKJJ8JpGzVqZB5//PHcVMa7v8Ya+l0/grivveDnT2AGCMo0DvJHxEqNon0TF9f/3XMOL32J0zBQnmEM2j/aHzuVYH9mPHTLBLgd5UKZJoEFZgxQAyaBBWZxcrLoNF0HtRi5jJ18k/LNN9+YXh0KfyINA+UZh4/+c0fkv+zj+pCSEyGjdYwDyjSIf/JgRL6xufLE/ClaND95N9sy/zOivXtHMTKNP73Mi6ax2T+py7oF7eMp2+ZPq4HydHnfXuYO6pGDeeI85Yu81o033ui9tgzvv/++dw5BdzrZj9Af7r33Xq8odKeJYq211jJfffWV9/qyrbLNKAsXyjQOd4wb5H3YonXViuv/rlz4Aq1jVCjPcr351F/Nio0qfwqictmfGUcd3AtuS7lQpklggRkD1IBJYIGJydGKHXbaHG5H2kiusr+YDPv27FHwE2kYKM84vPvvm+H6lyOuD6lLzjgWrmMcUKZBjukdfMqmTdZbs7ZNi+2zaZM3xb+M7gfPs1mMTCvzaIoI/1tyWSdZNzSNT7bN3tZSUJ6u+TM+8PqADEOGDIHLjUL+P8k3O/4g3ybaRezQoUNzzxgzderUxPaxkwOR/GH+j+/CLFwo0zjcPHYgXMdyxPV/99gy+5QWyrMccnaK3nviq76ljf2Zsf9++5of33kAblM5UKZJYIEZA9SASWCBicmHaNS/2CtJTsMig9yOH9oTbpMWyjMOcgT5ckUOBNGS/d4233xz78TF6Hmtv04cDdcxDijTIBOP7wXX0da3c/Y0VOcP2Qs+7+rbpZk587A94HOITCvzoOdcsg6yLrJO6HmbbJu9raWgPF2L5/7k9XXZp2/VVVeFy42DnFbIH+S0QjJODt6ZNWuWN072Y0PfbsZFrncup5SRYfHsH2AWLpRpHOQIcrm+P1pPrbj+744emN8FJE4oz3LIT83yGYfWOY3sz4wHbhoPt6kcKNMksMC0tG3V3HRo19p0zOjQtpVp3WIXOJ0LNWASWGDWFXTQQlp16NDBe7OQo1D7dNoRbpcWyjMO8hf+VpttBNe/0l56eDJcxzigTIPIVXOCfmYW8n9HTqZ/9uAe8HmXnE7GvUBAEJlWewoaWQdZl1IfprJNxa4uVAzK01WzOHs6nxdeeAEuNy7ys/dzzz3nLUt+TpQDie677z7vsRR+Qdcpj4v/LdPShXNgFi6UaRzkF52N1kmumC4HOrtCHFCeWnKgzI7blt7fOU3sz4wTDu8Dt6scKNMksMDMaN+mpRlyxGBz8YUTzJRJ15jrr51iJl9zlTnvnLPNgAMPMC13bQbn86EGTAILzLqO75PsB0ex07lEIefak0uALVq0yLTaqWmkExKjPONy9CGlv61L2kYbrOOdSgStXxxQpqUEnQzdt9GfVzej+neBzyErrqD/6bacaWUdZF3Qc7ZiJ3EPgvK0zZr2ROYjMXtqor///e9wuXHaeOONa8/fKP+//GHSpElw+ri9+GL20pVy1SGUhwtlGpde7fG16StJrgolp45D6xcVylNr4tnHw/WNywoJ7IZhf2Z06dAq8gUoUKZJ+MMXmG1btTBnnH6qV1T6heUVEy8z106e5D2+bspkM/TIwYFFJmrAJLDALHTP2YeWdTLhckhn7dZia28fIvR8VI888oj3YdS/f/+iV1vRQHnG5T8PXBP5p7aoTht2MFy3uKBMS+nZZlu4rq7110ruJ2Et7TrINqFtDYLytFW6wBSHHnqotzx/kJ/m119/fTht3F5/Xc71KefEnAfzcKFM43LNiP2993C0npVy8B7N4brFAeWp8fkr95R18YhySN4H9enm7TOOno/K/8wYMKC/eedfN8Pt00KZJuEPX2D277t/ppCc7BWT551zltl7zz3M7p07mH4H9DFXXj7RG3/NVVd6P5uj+QVqwCSwwCy0X8dMw4J1j0rOLSingJFvFuVqFGiaqEaNGuW9WVxxxRVmVJHrUmugPON04L76b+Hitt46a5ovX7sXrldcUKalDO8b7fyJaSTbhLY1CMrT5f9ELlfiQctNgv9TuQyaK/zEQb5h8s8dKfudoixcKNM4ddllS7iulbDmqo3NveccCtcrDihPjeMG7wfXN6q11ljN3DhxjPfNolx9DE0Tlf2Zcf0lo+D2aaFMk/CHLzCPP/Zor4gUB/TpVfDcSSOG1T7Xo9tuBc/ZUAMmgQVmnlyhJO6fr2Wb5VKTt542sHY5Fx5d+kjgMNq1a+e9WcgH756tmxZsWzlQnnH67L9/M002qnvNakSO0JXr9+61117mkEMO8Y6sPeaYY8zhhx9u9ttvP++ygNqDBuQAoyTPf+lDmZYyaUTwCdTrI9kmtK1BUJ6uxXNmeP1cLq249tqV2Ve6d+/e3jJlkL6Ipolbnz59ckuUc2F+DLNwoUzj9LezDjHrrqn7BjvO/7vyq0dS57/0oTxLefnRa02jMnYv0ZBtlUtNvv/MrbXLeeS2C+G0UdmfGYP77VmwbeVCmSbhD19gHtT/wNoi8sjDD6sd36r5zubMcad54+Xn8s4d2hbMZ0MNmAQWmHlB5yMMY/MN1vKORnf3h0yqwJQ36zlz5ni23XzjzHLD7auE8oybvDFvuB4uDtZZZx3vw0iumWvv91ZskCu5yNVBzj33XNOsWTOvn7mvKcXlVecNg+sSN5RpKQ9feGTmgyr951zVkm2RbULbGgTl6Zr/Q/7yjKNHj4bLj9vuu++eW6Lx7qNp4iR92N//UnYJmD39GZiFC2UaN/lDfO3VV4brncT/XSm4hh3QEa5LnFCepQzo3bXO+kaxY9PNzcO3TqizP2RSBab9mbHrTtua3z4Mvx8myjQJf/gCUw7wkZ/GpZCcMulqM+qk4eaIwYeas84Y5+1/KeNPOO4Y7oOZINSAQeQv80YxnVR9lZUamaH7tjEPFjkfpfZUM2HIX6IyyCXr5NyGaPmloDyTIH+hd2qTP9WNnMLk7rvv9r6ZsoeffvrJO2JYzkco+wyJRx991DzzzDPm008/LbhcX01NjXdU5D777FP7uuuvs5b5+w3nwnVIAspUY/vNKrNfXyXItqBtLAXl6Zr1yZOmZmn29D3SN+Sk5Ggd4lTpAtPe73Px7O9hDgjKNAnyi0yzLfOXjkzq/+5aqzU25x6xJ1yHuKE8g8gvMSutGM8J9ldfbRVzwdihZsa7D8Jl/fPG8+F8cfA/Mzp37mQ+fuEOuHwNlGkS/vAFpti9S0dz0YTxtd9k2saccrJp17oFnM+HGjAJLDCzTraOzm3btq0ZMGBA5i/n8n4ul+2TfZRuO/0guAzfaQd3g/PH4eqrr/beLEaMGBH6jRnlmRT5i/nSM4/z1l2O2J05c6b3QSMHN5x22mnetxpy7Vx3O32S+UYbbWSOOOII71uT+fPne9s/ePBg7/lee7Q3X7x6D1x2UlCmGn0S2v+3GmRb0DaWgvJE5s/40GtnGeRKOmgd4lTJAnPbbbc1v/32W3ZhNUvV314KlGlS5BeS4/bLnnEjif+77XfczDvoEi07CSjPINdedHLttoT9zJBvZ2Wf9A+fuw0uw3frVafB+eNgf2ZE+UMcZZqEP3yBuWf33c1lF1/kFZNyiqKLJlxgzj37TDPx0ktqv8E856wzvW860fwCNWASWGBm7dFyG28dt99++9od68u5SogceX7W4D1Upwc6at+28DXicOSRR3rrfsstt4Q+4hLlmaQn776sdv07d+5sdtlll4JtKof8RCdH0Utfk8cnHrE/XGaSUKYacmCWuz1xkkzkA1D4+SQl7EFmKE9o2uNmyYLfvb4uw5lnngnXIy6VKjDXXXdd7wTu/iBXLYLbXwTKNEmXWRcJiPv/7v6dol/2thwozyCH9M1eyCDsZ4Ycef63a89SnR5owmlHwdeIg/2ZEeUMGyjTJPyhC0w5kbq/n6UUl4cdfFDtT+FtW7cwJ48cUVtkHjXkiDrz+1ADJoEFZtZ2m67nreOll17q/WeT4ZRTTqmzDcgGa6/mXWYPvS7SvcXW8HXisOuuu3rr/r///c+03m4TuPxSUJ5JGjfiULgtcdhpuy3gMpOEMtW4+Jj8T4PlkG+Jtt56a7Pvvvt630Jcfvnl5p577vF+hnz33XfN119/7X0jNm/ePO8nTCH3ZZw8J9PItDKPzCuvIa8lrxn0DVQQ2Ra0jaWgPIuZ/fmzpmbJIq+/yyDfmqF1iUMlCswNNtjAvPnmm7mlGLPo92/gdgdBmSbp0B4t4LbEQS52gZaZFJRnkDbNt/PWM8xnxuabbGDeePIv8HWRQft3h68TB/szY6/dW8Pla6BMk/CHLjDlwJ2rr7rCKyAnjD/PtGpeeOUeOWXRpKuv8p4/4/Sx3oE/9vM+1IBJYIGZJQfkyDo+9thj3n822U9o5ZXxjuw22d/yhlP0xaX8rLR+piBFrxUH2Wlb/pqWnbY332i9UAf6oDyT1KFVcj8Ny8E90168Ey43KShTDXkja9wof83rYrbaaivvZ8Rrr73WvPLKK7XfniQxyGvLMmRZskxZNlonm2xD2DdllGeQOV+95P2M7A9XXnllwXXDtdZYYw3Tpk0b72fOk08+2UycONE7HdE///lP8+CDD3ofvv7w/PPPm9tuu837aXHs2LHe/pLy7d2GG24IX1tj5513Nl999VVuCcYsnvOj9y0t2uYgbp5J23GL/H6YcZOfj+8842C43CSgPIPIATmynuV+Zsj+lq8/cQN8TUR2I9qsSXL7Z9ufGU233jz0gT4o0yT8oQvMju3amCsmXuoVkJdfdqm3L6b9/MD+fWtPuJ6WAlP2lRk/fnyievTokeoC03+jlB2e5S9S7YfU8L7lHd0oJytGrxMn/1uQFi2am7vPOgSuRxCUZ1K+eeMfZsWAoqpx48amZcuW5uCDDzZjxozx+tKFF17o/SQqpzzZY489Sp70+qbLT4XLTgrKVOuQPep+IyTFj/x0eNNNN5kvv/zSa9ugQfaD+/HHH81bb71l/vWvf3lFkhREN9xwg5kyZYpH7ss4eU6mkWllHpm31CDrIOsi6yTr5q6vbAPaNg2UZylzv36l9qAfGeSclVtsUfyyfXL6nNatW5tTTz3VPPDAA+aLL74oONgkyiAHtfzf//2f10/33HNPVcEhP1HOnj079wrGLJKDekIUlwJlmpR/nDfYrBBwYGQc/3dPHZTMdccRlGcQ/w/jcj8zrj5/OHy9YuTiFOh14uR/ZrRs2cJMf/luuB6loEyTIAVm5WqWlBWY8nP4qJNGeAWkuOD8c82gAf2882HKKYvkij7+c4MPGVRnfh9qwLjJ5fI22Wg98+9//9vrXEkOM2bM8N7Y5aoHaF3ihhowSN/O2aOZ5Q3R/c9XzKbrreldtxy9XjF9u+SPmk7Krbfe6mUu3zhdcuy+cD2CoDyTgk4g3KRJE+/0M/JNkb/jf9AgxcGHH37onSxYdrZ39y+Men63cqFMteQyeB12yn4zIn1x6tSp3qlc0LBkyRLz3nvvmdtvv90rluRcjXKAiJyg297+csi88hryWvKad9xxh7cMWRYaZN1kHf3/N7LuUS7lh/LUmP3F82bpovw3ubNmzTInnXRS7Ye+3Pbq1cvbnp9//jk3FR5km3744Qdv1wHpg08++WSBp59+unbXg1LfHsvzko8UkW4xLge43H///bkps8PC377IFJdT4TZqoEyTgi4YEff/3Sjn8y0XyjPI8CF9vXUs5zNju603NT+//xB8vWJGDM0uJ0n2Z8bUOy+B61EKyjRu8t6y3lqrVrBmWa5iB5q5NWDRg3zkZ/Lzzz27tpAU/n6XvpNHDDNtWu4K5xeoAeMkOxb7VyAYOnSoef/99xN12WXZAzn27tbW/PLBw3Cd4oQaMMjkkQeY5co8AnDcod3haxVz3/mDE7sMpe3000/3/oNccMEF5oQ+HeC6BEF5JkUOwvHXW96o5fJ/cm1cf5Bv1L7//nvvQ/3GG2/0+tHFF1/sfQsnP11+9NFHZvHi/LdXMr38nDlo0CDvDxp53U03Xj/ydXbLgTIth/zRIudklW/C7EG2U86NeP7553vf/qy+eunrgcdFliXLlGXLOtiZyyDrKutc7h9cLpSn1qxPnjKLZn2XW6Ps8MEHH3g/m3/77be5MflBCkk54ln6knyj1rVrV69AKucndtlHVQ7MkeJITiAu32TJh5/83OgOMu4vf/mL9+3LyJEjC84TKd/AzvvuTbhd5UCZJkUOwvFzSOr/rlyWVHPgZBxQnkFefGiyWb7MfZTvuGYcfK1ivnvzvsQuQ2mzPzMuP+cEuC6loEzjJP3Av9JeJWuWtttvGuqcvuVya8CiBaaQ4nFAv77mtFNHm0svvtC7ROSE8eebk08abvbt2SPwHJgCNWCcLjz96IIOVklDBu2T+Ac+asBSDizj28Wmm6xb9v6Nx/RK5hrkrr59+3pvFvKGH+Z0MSjPpMhBOFtuuaX5xz/+UfszpXxbJj/bHnfccd6BJu63Gi65msv+++/v/RX+++/5I4vlmzc5p57M/7+n/gqXnwSUabnkL/XJF55hpk+f7mUjPzNW6qo1GrIusk6ybrKOUy46I9I3lz6UZ7nmffdG7eUk3UEKzUmTJnn9YrXVktsXulGjRt5+mfJTm3xDFzTIZSDLORVREJRpUuQgnOT/7y5j/jq6P1x+3FCepYw86kC4XUjLnZuWvX/jReOOga8VN/sz4/jBfeC6lIIyjdPRvZI7+0op+7TdLvE/dNwaMLDAjAo1YFxuu/p07+AHFGSlnDf6SLhucUENWIp8QA7sukvJy0XKm974oT3haxQj+0KuXoFvL8VOO+3kvVm8/fbboY4kR3kmQfa/XGH55b2reMggRzfLtxvywYS2S0OKhmHDhplvvvnGe035RkS+kfrrxNFwHZKAMg1DrrtciW+8o4rzGtEozzCyJ2PP/qwv35LJN2ayT2TYo+KjkCJLLoso+73aP6lLETzv+7cz6xv+J3EXyjQJsv+lvE9W4v/u6IGV2Q8T5VmK7GZ2ynEDS14uUvrAAzeNh69RjOwL+ee1KvMrhf2ZEfZIcpRpXE4/pJt30Bda90o5cu/WcN3i4taA9bLAlHMONl4pnqsPRCGdJcmDL1ADav11TH8zqHtz70S/W2705zrr3nwbuQwjnheRbzrleuTu6yRFfs6U/Z/kNDRbbrweXKcgKM+kyP4+3Tq19H56lfPJoe0JQz6s5MOvS8c25opzTyh7v6coUKZhjT04eym6HXbYwduPT86zlwayLrJOsm6yjmjdw0B5hlWzNPtz7UMPPVTQN5A///nPpn379uaggw7yDkiRn9Vlf035dk5+/v/Pf/7jefbZZ819993nndLpmmuu8Q5YkROFy6mL5Of1Ut/Y2ae0mfPFf+B6R4EyTYrs391y200y/3fPS+T/bpvmO5kT9u8QebcLLZSn1ptP/dWMPXGQd2GHZttvWWebunZsXtavdvJNp1yP3H2dpNifGTtuuyVcp1JQpnGQc62m4TK68n87yYPO3Bqw3hWYct6tSuzPoSVHDz92x8VwXaNCDRjGlJP6et9Y+uu89morm1vGDoTTFjNknzYF210Jn3/+ufchtvWWm5sHxuNLVhaD8kzaCw9OMkMH7WvWXjP6z5byreieu7U2d046o6KFpQ9lGkWvTrsUHGWclkHWSdYNrXNYKM+w/AJTvr0s6B8rrOAVk3LeTCk+5RuzuI4ilwOIZJ9DOVq6Z8+eZtVVVy1Ytl1gzv78ObjeUaBMkzZpxP5m33bbm9VWXrFgW8OQb0VbZ4rWMw7tXrHC0ofyDOOlR6YU/KGxwbprm/eeuQVOW8z5Y/QnbI+L/5nRdJutzQ9vPwDXKwjKNCo5v3SafsWRsyaEPcdvKW4NWK8KzE9fusvst++e3g7U8he37CR79NFHm2OPPdYcf/zx5sQTT/R+nnANHz7c2yFdQ6ZFryGvLcuQZcnO9LJs+QbkkEMOMb326Wleeew6uM5RoAYMQ7593Kv1tqbxiiuYlk2blHVCdSHf7lTjq305cbYMcn3ZUpeudKE8K0WuxSt/dMjJ16VI3HC9tUt+K7TqKo1N61238w5ak0uqyTWC0WtXCso0iuP27+Tt55i2QdZJ1g2tc1goz7DsAlP2idxvv/3MXXfdVfIocjkJveyrKT8Xyv8j2afQJgfxvPHGG94HcqnCX74VkqPI5T1vzTXXbJAFpu/BC47wPnzl5OtSJK69+soFf5wj8r4qF7mQgzfkErp/C3FatbigPMOQbx8P77+X9760R+eWZZ1QXdxy5diq7MKW/8zoXPLSlQjKNIq7zjw48xnQIXU1S88e3cx1ow6E6xyFWwPWmwJT9hPp0m5X79QdaRvkyMF9e3aP/XrRqAGjCPPX9IVH720aBZwnLkl33nmnl6+cq3Di8b3g+hWD8qwW+VlJCkbZtWON1Vcp2EbZAf7df99ckbMSlANlGsXuu27lnQxZTsYtl+JLA1kXWSdZN7TOYaE8w/ILTCkW5bRD7iBHkb/88stm8uTJ5qijjjKdOnXyTh3kH8GsIZfdlEscynk15aCnSy65xPsG0z5gxR/kKHJ//0IZGlqB6ZLdiKRglJ84V2lcuFuWHPB489iBFTk6VwvlGcVP75X/68kjt11oVlqxOruw2Z8ZT90zEa5fEJRpWHI8xK5NN01tzdK9S/vYT1/k1oD1psD88Z0HzIqZv+DlxMqvvfaad1JlOQxfrnkr30LIFSTknG7fffedd1oJOeGynDBY/tIXcjoNm+ynIdzx/vRCXkNeS15TXluWIX/xT5s2zTt1iHw7IKcIeeKJJ7y/7OUnUrTuYaEGrCQ57dGqjaP/ZBTWRRdd5P1nkEuXyQ7SaB2LQXlW04fP327aNq+7j9eaq69a9o7zlYAyDevv5xxm1l2z8GfWNJF1+/u5h8F1DwPlGZZfYNqDvBdJQYl+vo6T/AzfoUMHb99iOSJaPpTcoaEXmOL2cYPM9putXycfeW8s90DJpKE8K0lOeyTvaW5WlWJ/Ztx+zelwHYOgTMN64IIjvAOn0lyzyK4haN3DcmvAelVgyn5pqFMJ+QmyEtCyfXK1ArTuYaEGrBT5SVpOBou2s1Lk630Z5NrSR+3bFq5nMSjPapCrPl18xjFmrTWK75cpux/IidTf+dfN8DWqAWUahhRu22+xkXeORbkqCtr+apJ1knWTbxri2l8O5RmWX2DKqXPkwBw5j2c1jiIXchS5FLb2+TEbcoEpVz85pne7wP0y5TNBTqR+86kD4GtUGsqzUuQnabnoCcqpUuzPjAmnHQXXMwjKNCwpMIPO5uLWFklBy/bJVfnQuofl1oANpsBMg4ZSYMrpO7bauO6R55Um+5vJcO+995r+u5d3IAbKMyz5iVt2GJdTbsibqOzsLsXgW/93o3duSrkm72uP3+Dthys7x//fPZebGy49xRzSd4+y/pqXEx5369TCK0jlZyb5NuDlR6/1XluWIct6M0OWK8t//5lbvWuUy6mS4v6JHWUaxm67bOXtvyeDFCayL6F8CDRt2rTkm18SZJmybFkHWRe/WJJ1lJ880TaUC+UZll9gPvzww3B7bOutt5534M9hhx3mHfwjV5aR/TUfeeQRb980m3yD8be//c0rGM8++2xvv7Bu3bqZTTbZxPvJHL2+rz7tgyk/ccsBgnKKNfmjWQ5ulGLwxjH9vXNT3nBKv4wDvf3R5GDIy0/obU4ZsJvZo+U2Zf16Ixe4aLHNxl5BKrsVya8/157c13ttWYYsS87sIcuV5d962kDvGuXyXhvnT+woz0qQ96Bddix9jf+k2Z8ZJx/TH65rEJRpWKUKzDRggZlTHwrM5++v/wWmvNnJzu1o+ypN9gmTQS7Z1qNVeZdbQ3mWQ/aLvPTM40zPrm3MRuv/2Sv+tH8VVoq/LvIN6OqrreJdV/jUEwaZf//jyrJPhuxCmZZLPmTlAAl/x3t3kJ9x5Fu5sWPHeud33GCD7LX04ySvKa8ty5Brlssy0SDruO0m68LtKBfKMyy/wHRPU+SfBH3cuHHm0Ucf9X4WQz9hhxnkZzg5lZHsi7nvvvvWudpS2gtM2S/yuP3amzbbb2r+vPrKXvEn/dBnb0u15NfnT2aVlRqZHbfYwDut3JUn7ucdlIm2SwPlmTT541YOZkTbWWn2Z8ahB/aA6xsEZRpWvSgwh7PA9LDArAw5ESvatmrYaqutvDcLuYpIux02g+tbDMqzFHmjlP12OrVplvhR80kXqVtttpE595QjQl83H2VaLvnAlHWR61fLN2TyLZz98yoaZJ+iV155xfsGYuLEid41oeXoS7lSivw8LAextGvXziP3ZZw8J9PItDKPzCuvIa8VNMjR07JOsm5SRK21WmO4HeVCeYZlF5hyjfUDDzzQ3H333WbmzJne+GKDHEUu+17J/lbPPfec942lnA9TrnIi32jKuJdeesl8+umnXpsEFadyAnK5frkcjbrWWmulssCUP4xlP+1mW26Q+P+tpIvUjdZZ3RzRs1WoAzBQnkk7b8yRcDuqwf7M2Ld7O7i+QVCmYbHArIcFpuxwLm+W/hukHEH56quvem+kctWEN998E5KdW995552S0LxCXluWIcuSDy9Ztpy0+KmnnvKuUStv/vW9wLxj3CDvlBuoI1aDXB9ZrmAiR9DusPkGcJ2LQXkWIz+B3zn5TLPtVsl/c9t0yybeaYjkgLB9urVNvJBdbdWVzWnDDvb2BUXbXgzKtBxyVZx11ig8Yl6suOKKZrfddjPnnHOOd/LvUoVSnIMsS5Ypy5Z1kHWx101OhBzHJf1QnmH5Babs/C878LuDFJL//e9/vROmy1HkclCOfGtbzn6aUpDJ5Q7lWtxyFLkcKFGsbeQqPnLwgD9Uu8CUn8DPPGwPs8l6a8Jti1OTddf0TkMkB0a03WHTxAvZlTPvxQfv0dzbFxRtO4LyTNJH/7nDO5URWv9qsD8z2rXYAa5zEJRpWH6Bmeaa5Q9dYE6+cKQ54fA+nmMP621WXrmxd1qONA4tWrQw/XvvXru+Z448DG5TOVADJumwPVvC/7TVIv8B5BQPYptNkykwZR9G+RkcLT8uq2T6be8e7c1dU86ss6+k7Gcp577ceMN14bxx2WLTDc2jt19UsOwgKNNyHL5XK2+5cnWZoGJH9vfbdtttzYABA8x5553nXV1GjricMWNGqBOHyzwyr7yGvJa8pry2LCNo30JZR1nXTs22gNtTDpRnWH6BaQ9ffvmlueqqq7yf/ldeeWW4PXGQUx3JAVCyj6YcAZu2o8hlH0b5GRyte1waN1rBuxqaFLHuvpKyC4ic+3Jd8IdUnDb88+rmoqN1J8ZGeSZJPufQOleL/Zmxy47bwHUOgjItx8h+nU2fTjt6enfYwTuIMM01i5yizV9f+fxH21QOtwZMdYEpH8puB5KfxOQEoqNGjTKnnnqqtzP7GWec4X0rIZfmGj9+vLngggu8q1DIPkRCftKRn85scpSZcMfLtP588hoTJkzwXlM+qGQZclk1WaYsW06FICc0lQ8w96/ZzTfZAG5TOVADJkW+CUCXlKw2+dZGioZtt2jirSNadwTl6ZLicqMN1oHLDSJtLd+myzV2N2uyvtmx6eamTfPtzO4ddvX67GEH7mlOOqqfueys48wTf7tUdUUJ2Wfy1anXm+suHuVdrm3IoH1M3326mO6dWnj7Vsql27bcbCOz/jprZd60Vgz1zaec+Fh71SmUaTm6Nt/aHHfccV5RIvs9Tpo0yTuIRE59g9YNkW8Y5aATOXq5a9eupnfv3qZfv37epRCF3Jdx8pxMI9O630oGkXWRdZJ1k3WUdR0zaiTcnnKgPMOqWTw/93GQHR577DHv20a0PUmSfT7l0pPuMHv6M3C9o0CZuqS4RN+QlyI/b8u3SquvspJZf+3VzOYbrOWdJH3XrTfyCsk9WzU1/Xbb2duH89LjeqmuICb7TF4/6kAzqn8Xb7eQfdpuZ7rsvKVp0bSJt2+lvK9ulCkSZReMFVdYPtQ3n/L//eJj9oXLt6E8kyK//KBLSlab/5mx847blnVpS4EyLYf0IXd96kvNskHm/wPapnK4NWC9KzDri/pWYMpPmmncX0TO3SUf/Ltk3izKOY0MyhORy5mVesNfb501zUF9upmrzhvmFYxyJLlcrSfqgTRhyBumfAv69et/944wl5/bjx/cx2yTKcDRutukWNVePg1lWg7Zl1cKN3eQn13lYBt5w23WTPZ1rVyfk2XJMmXZsg7oJ+B777wFbk85UJ5hzf3mVbN00bzc2mUH2Wfy1ltv9c6DWU5BXS7Jq02bNt6HmHtwVM3SxWb+j+/BdY4KZYrI5WtL7Q+55qqNTbcWW5thB3T0CkY5klyu1hPlQJqw5A9k+RZUTt0lR5jLz+19Ou5omqxb+tLHUqxqil2UZ1K+fO3eVB4X4X9mtG6xS9mX2UWZlgMVmPUFC8x6pL4VmLJfUdI7r4ch+63I0LFdm7KuR47yLOaaC0ZkiuvCn3Gl6JRvJP/xl3NjPwVQEqTwfO7+q73Lu6GraOzfs5O3HzOaF0GZlkNOv7LtFht7R2/LvkDo51UZpMiTq8ZcdtllZvDgwd5RoHIgibv+5ZLXkNeS15TXlmWgglIGWTdZR1nXYw/oArenHCjPSKY9YebP+MAsdb7NlEGutiNHkY8ZM8b7JjfKt5tyVSPJ7IQTTvBOYYSOuK9ZusQs/HW6mfXZ03hdY4AyLWbEgZ28o8Tt7ZD3MflG8twj94z1FEBJkcLz6uF9vMv5oqumyW4bsj8fmteF8kyK7Ece5tvYpPmfGV06dyz7euQo03KwwCysAVlgJqS+FZiXHrsv3I5qk9PYyNChXVtz3/mD4bojKM8gd046wzReKVuYycE+96fw6jpacn5M2R/Yf/M/YmDPsotklGm55AooclSvrMMWW2zhXTNXfuItde1rKfjkCHDZyV2OXpZzOU6ZMsX7CUh+9jnrrLM8cl/GyXMyjUwr88i8xQpaf5B1kHWRn4tk3WQd5cMhjpOtozxjMe1xM++7N83iuT9ltqD49skBDi+88IJ3tLn8rC0HGfjXLBYjRozw9quU7G6//Xbv2uRyxLmczL3YsGTB716RO+uTJ/G6xQhlGuSMQ7t7B2hJG8rBPuOH7AWnqw/k/JiyX5z/x37PNtuVVSSjPJPy+F2XeuuYNv5nRqeOHcx3b94H170YlGk5WGAW1oAsMBNS3wpMOcEw2o5q69ixo7c/yYorNvK+FUPrjqA8S5ETpJ8z6nDv52/0fH1zz3Vnm3EjDi17PySBMg1Dvp254sT9vP3aNlt/Le+DU/bnk6OdZZ+g+++/3ztopVRBGGWQ15ZlyLJkmbJsWQdZF1knWTdZx3L28Q2C8oybfIM474e3zaLZ35uaJfEfRFBTs8QrZOfP+DCRA3mCoExLkfcvObBMfv5Gz9c3Zx/ewxzao0XZfRLlmRR5v0Tv2dXmf2astNKK3gng0boXgzItBwvMwhow1QWmfAUv12muj2RfPbRN5UANmBT5tkmuupJmaT5dR0ODMo2DfEMjR1rKfnFykIX/TY38tCvntRw6dKi3o/qdd97pnfxczmcnp+iRIzFRESrj5Dk5clymlXlkXnkNeS15Tf9nY1mWLFOWfVJmHWRd0DpGhfJMmhSB8777n1nwy6dm0azvvG8ca5YskIBySYEh81zNkkVm6cLZZvGcGd5P3/N+eMfM+fIF8/u0qXA5lYAyJR2UZ1I+fP5206/XbqlW6dOzya5mcn36+kj2UUbbVA63Bkx1gflHhxqQdFCepIcyTcJdZx5szjtyL+/bp67NtzLbNFkHXvtZfu6XU37ISdvldEJC7ss4tB+YvIa8lrymvLYsQ5aF1iFuKM9qmvXp/0HVLCKDoExJB+VJeihT0nNrQBaYKYYakHRQnqSHMq2k+84b7F3HWU7NMu7Q7mbkgZ296zzL0emD92zpkfsyTp6TaWRamUfmRa9ZKShP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oCJFphoBUgP/QcgPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BrwD1Ng3nnGwWb0wN1Mn447mk7NtjAtmjYxnXfewvTbbWdz9uE9zH3nD4bzVRNqwGqZ9uKd5i+XjTbHD+5j+uzVyXTv1MIcsHdnc9LR/cw9151tvnvzPjhfNaFMq4F9Lxr2vfDY96Jh3wuPfS+a+tj33BqwwReYU07q63Xu5Zdb1iyzzDJFrdK4kendYQfvPwV6nWpADVhpLz0yxezfs5NptMLyMDffGquvYo49rLf3nwK9TjWgTCuJfS8a9r3w2PeiYd8Lj30vmvrc99wasMEWmI9cOMQM7LZrbSf/05/yDSP3Xf5z0ulPGbAbfM1KQw1YKb9+8IgZffxAs8Ly2U7+pz/9ycrvT3X4z0mnv+HSU+BrVhrKtBLY96Jh3wuPfS8a9r3w2PeiaQh9z60BG2SB+cD4I0zb7Te1GiffmYPu+4/lVv6jPHoRfv1KQQ1YCT+8/YDZu1tbK5vCjl7svv9YbuU/ysyPHoWvXyko06Sx70XDvhce+1407Hvhse9F01D6nlsDNsgCs8suW1qNkL+179vP28/ZjunVDr5+paAGrIQD9+1Sm4Hdge379vP2c7aLxh0DX79SUKZJY9+Lhn0vPPa9aNj3wmPfi6ah9D23BmxwBeawAzrWhu12brdjF7v178tX/VcN6wOXUwmoAZN21XnDrAwKO7fbsYvd+vflq/5n/3kVXE4loEyTxL4XDfteeOx70bDvhce+F01D6ntuDdigCsy/n3OYWWOVlXJhZ+XDz9+3ny813Q6brQ+XVQmoAZP01Wt/N+usvUYuh3yn9h/79+3nS03XrsUOcFmVgDJNCvteNOx74bHvRcO+Fx77XjQNre+5NWCDKjCP7d3OCj3Lv++Pt5+379vT2vfl9vITesPlJQ01YJIuOeNYK5N8J3Y7sDvOnda+L7dP33s5XF7SUKZJYd+Lhn0vPPa9aNj3wmPfi6ah9T23BmxQBab85eN30GzY+Vt0Hz2Hxu3faSe4vKShBkyS/OXjd9DstuMO7E5jP4fGnXjE/nB5SUOZJoV9Lxr2vfDY96Jh3wuPfS+ahtb33BqwwRSYD1xwhGm0/HKZcOt2XLn1yWNfscf2tHLbdJN14TKThhowKT++84BZacVGmW2u23H9PPzHvmKP7WnltuXOTeEyk4YyTQL7XjTse+Gx70XDvhce+140DbHvuTVggykw/zqmfy5gzH7OvV/sOd+aqzaGy0waasCkvPnUX3Pbnu+8Nvs5936x53zr/nlNuMykoUyTwL4XDfteeOx70bDvhce+F01D7HtuDdhgCsxrT+5rBV946993x/vj0GObnAgWLTNpqAGT8t9Hr7Wyyndae5w73h+HHtvkRLBomUlDmSaBfS8a9r3w2PeiYd8Lj30vmobY99wasMEUmLeMHZgLPE8e++P8+/Zj+9YdZ1trtYb/19R7z9yS2/58J/W3375vP7Zv3XG29ddZCy4zaSjTJLDvRcO+Fx77XjTse+Gx70XTEPueWwM2mALz4QuPNCuvuEImbLtR8vzH9q09jf/YHSe3zbbcAC4zaagBk/LLBw+b1VZdObO9+c7qd2K3I6Np/MfuOLnt1KYZXGbSUKZJYN+Lhn0vPPa9aNj3wmPfi6Yh9j23BmwwBaZotW2TXMD5jure9x+j6RB5/tAeLeDykoYaMEk9urTK5ZHvqO59/zGaDpHnx404FC4vaSjTpLDvRcO+Fx77XjTse+Gx70XT0PqeWwM2qALz1EG7ZwKW8POyjZG9ddnT2OPs+8su+ydz45j+cHlJQw2YpJsuPzWzzXU7q3/rsqexx9n3l1tuWfPW/90Il5c0lGlS2PeiYd8Lj30vGva98Nj3omlofc+tARtUgfnQhCPNJuutmQu6UL4Bij92x8vtbrtsBZdVCagBk/Tz+w+ZbbfaJLf9dTu9PR49dsfLbb9eu8FlVQLKNCnse9Gw74XHvhcN+1547HvRNLS+59aADarAFBcfs49ZbtllrdDzt+h+seeEXALrttMPgsupBNSASXvsjovN8sstZ2WT78jofrHnhFwC68PnboPLqQSUaZLY96Jh3wuPfS8a9r3w2PeiaUh9z60BG1yBKYbu2yYTtgSf78D5hil+a1th+eXMhKP2hq9fKagBK+GCsUMzGRR2YLm176Nb24qNVjAP3TIBvn6loEyTxr4XDfteeOx70bDvhce+F01D6XtuDdggC0wxZB/p8BK8NES2obKNgvnPyW3jFVcw5xzeA75uJaEGrJTzxwzx9oXxO28+v/w4m/+c3K66SmNz7/XnwNetJJRpJbDvRcO+Fx77XjTse+Gx70XTEPqeWwM22AJTjB+yl3c+LbtD2+xx/v0tN/qzuX7UgfD1Kg01YCXdf9N473xadoe22eP8+82239K8OvV6+HqVhjKtFPa9aNj3wmPfi4Z9Lzz2vWjqe99za8AGXWCKNttvmmuMPP+xPd6/P3jPlvB1qgE1YKX17Noml022w/ud2r6175910mD4OtWAMq0k9r1o2PfCY9+Lhn0vPPa9aOpz33NrwAZfYO6y1UaZRsh25myDZPn33XF9uzSDr1MNqAErrUu7XTLZZDtzNqvgDj9iaF/4OtWAMq0k9r1o2PfCY9+Lhn0vPPa9aOpz33NrwAZXYN53/mBzfJ/2psU2G5t11lil9ug2v0PbHRzdyo7G66+9munUbAtz+iHdvKsVoOVUAmrApH335n1m4tnHm26dWpiNNlin9ug2v0PbHRzdyo7GmzVZ3/TZq5O57erTvasVoOVUAso0Sex70bDvhce+Fw37Xnjse9E0pL7n1oANqsCceHwvs26mg0voPtSp0Tj7Of+xaNpkXe+aq2h5SUMNmKSn7ploNt5w3dptz2ZSt1OjcfZz/mPRollT75qraHlJQ5kmhX0vGva98Nj3omHfC499L5qG1vfcGrDBFJhy5v9VVmqUC70uf7zfCL5iz9njN11vTXP/+MPhcpOEGjApcub/1VfLvlHYndbuvP6trdhz9vjttt7U/PDW/XC5SUKZJoF9Lxr2vfDY96Jh3wuPfS+ahtj33BqwwRSYvdrvkAs3Lx98/rH7vPZ2VP8ucLlJQg2YlKMP6ZXb3sIObo9Dz2tvr7t4FFxuklCmSWDfi4Z9Lzz2vWjY98Jj34umIfY9twYsWmC22KWZOerIw83YMacEOnnkcNOm5a7wNVADJmXXrfM7Fvu3/n17vKvYeGG/xoCuu8DlJgk1YFJ2a79rZjsLO6h/3x7vKjZe2K8x6tgBcLlJQpkmgX0vGva98Nj3omHfC499L5qG2PfcGrBogdmq+S7mrDPGmeuvnRJo0tVXmfZtWsLXQA2YlAM675QLtpA7Lt8Ahc+h6ez7Yw/uCpebJNSASRl25AG5ba7bYd3H/jj7OTSdff+WK8fC5SYJZZoE9r1o2PfCY9+Lhn0vPPa9aBpi33NrwMBvMA89+CAz/MTj65BvLaWwlALziomXmXatW8DXQA2YFLl+qVzH1O6ocutzO7A7nX9rT+M/3qbJOubBC46Ay00SasCkyPVL5Tqmdkf1t99+7Hdgdzr/1p7Gf9x8p23MjHcfhMtNEso0Cex70bDvhce+Fw37Xnjse9E0xL7n1oCh9sEcNLCfuXbKJK/APOaoIzPF6E5wOtSASZo88gDTZF1pMD/0PPdxsfF+A/n3m2+zsbnrzIPh8pKGGjBJLz402WyzRZPMthfv2C40nT9Obrt2bG4+efEuuLykoUyTwr4XDfteeOx70bDvhce+F01D63tuDVh2gSk/h190wXivuLz8sktNp/Zt4XQCNWDS5BxaYw7a3bv8VDb0PP9xvkEKH9vjWm+3iXfh/UcvwsupBNSASZNzaN04cYx3+alsHnU7dj6rwg5uj9tr99behfdnfvQoXE4loEyTxL4XDfteeOx70bDvhce+F01D6ntuDVh2gXn4YYeY66ZM9grMIYcPhtP4UANWwqMXDTFbZTq725Fddme3b8VerbeFr11JqAEr4bcPHzU777BVJofCjuyyO7t9Kw7vvxd87UpCmSaNfS8a9r3w2PeiYd8Lj30vmobS99wasKwCs1OHtuaSiy70istLL77IdGzXGk7nQw1YCRcevXcu+EL2OPd5/7HcipUaLV+1r+l9qAEr4ZHbLszlke24Pnuc+7z/WG7Fyo1XqtrX9D6UadLY96Jh3wuPfS8a9r3w2PeiaSh9z60ByyowZX9LKS7F4EMHwWlsqAErYactNqgNvVhntu/bj+3p5Sg59PqVghqwEjq2zh4dmM0Dd2b7vv3Ynl6OkkOvXyko06Sx70XDvhce+1407Hvhse9F01D6nlsDqgvM3Tt38Pa5lOLyognjTYe2reB0NtSASZNTG2RDzzeE/xh1aHec/bjR8suZG045EC6nElADJk1ObZDd/rqdGXVod5z9eKUVG5nXHr8BLqcSUKZJYt+Lhn0vPPa9aNj3wmPfi6Yh9T23BlQVmHKUuJyeyP/28uCB/eF0LtSASbrzjIPNWqs19sLOBo7Zz/nTonnk8Xabrle1i++jBkzStBfvNOuvs5aVRb4D2+zn/GnRPPK4TfPtqnbxfZRpUtj3omHfC499Lxr2vfDY96JpaH3PrQFVBWaPbrubq6+8wisux593TtHzXrpQAyZFOmSLbTbOBV5XvjHyj+3n7XH2tHLbf/fKX1FAoAZMinTIbp1a5LY732Htjms/h6bzx9nTyu3Jx/SHy0wayjQJ7HvRsO+Fx74XDfteeOx70TTEvufWgCULzJa7NjOnnDzSKy7l6PEBB/aF0yGoAZMgpzXQXBfVH+c+9se50+fv/8mc1K8zXHaSUAMmQU5roLkuqj/OfeyPc6f37y+77J/MlAtPgstOEso0bux70bDvhce+Fw37Xnjse9E01L7n1oAlC8y99+pRe9Wec88+y7Rt1RxOh6AGjJt09H677VwbdDbguvf9Duw+h8bZz/n3l19uWXP6Id3gOiQFNWDcpKOfdFS/2u3Pbm/dTux3YPc5NM5+zr+/wvLLm9uuPh2uQ1JQpnFi34uGfS889r1o2PfCY9+LpiH3PbcGLFlgHjJogDnt1NGe3vv2hNMUgxowTnLurd4d8n9FFbv12Y9L3Zdbd/xyyy5rRg3YDa5LElADxknOvXXsYb1z25nvmO6tz35c6r7cuuOXX245c/0lo+C6JAFlGhf2vWjY98Jj34uGfS889r1oGnrfc2tA1T6YYaEGjIvs/9G95Ta5QOt2THTffiy3Pnc6+779OHv7J3NM73ZwneKGGjAusv/HwQd0r90m/zbovv1Ybn3udPZ9+7Hcylf3F59xDFynuKFM48C+Fw37Xnjse9Gw74XHvhfNH6HvuTVgvSwwH5pwpOnUbItciIWdUzuu2Hh7nDu9Pf6QPVrAdYsTasA4/PTeQ6bPXp1y24c7aqlxxcbb49zp7fGnDz8ErlucUKZRse9Fw74XHvteNOx74bHvRfNH6XtuDVjvCkzZ/8P9K8q+b99qxhV73n5sP2+PP75Pe7iOcUENGJXs/+H+FWXft28144rNYz+2n7fHTzz7eLiOcUGZRsG+Fw37Xnjse9Gw74XHvhfNH6nvuTVgvSswzx7cIxNU3c5X6jYImidofn9coxWWMzePHQjXMw6oAaO6+7qzM+tet/OVug2C5gma3x/XeKVG5t1/3wzXMw4o0yjY96Jh3wuPfS8a9r3w2Pei+SP1PbcGrHcFZvsdN8uFVdgp7U7ojrefR+P95+xbNE5u3ecP36sVXM84oAaMqneP9rltKOyUdid0x9vPo/H+c/YtGie37vPnjDocrmccUKZRsO9Fw74XHvteNOx74bHvRfNH6ntuDZjaAvOGU/p5X4fLEWt7td621pqrNs4ElQ0tG1ye/9h/zn3sTutOY9/a07m3Pnm8yXprFqxf387NzMn9u8Ry0X7UgFqvP3GD93W4HLF2eP+9aq23zpqZ9a7b8fxx9nPuY3dadxr71p7OvfXJ42232qRg/YYP6WuuvejkWC7ajzLVYN9j30PbVQ6UqQb7Hvse2q5yoEw12PfY99B2lcOtAVNXYN4xbpD3F5MbjM3viL6g8eixPz1iT+s/du/709jPueSaqn067WgeGH8E3E4N1IClfPSfO0yvPdp7R46h9RKSrS1oPHrsT4/Y0/qP3fv+NPZzLrmm6gmH9zE/vP0A3E4NlGkQ9r08lGcp7Ht5KNMg7Ht5KM9S2PfyUKZB2PfyUJ6lsO/luTVgqgpM6ejrrbWqt7F2hwpiT4vuy637esXGoefQffcWkedEsy038I7AQ9tbCmrAINLRN9lovdx65TtUEHtadF9u3dcrNg49h+67t4g8Jzq1aeYdgYe2txSUaTHse4VQnkHY9wqhTIth3yuE8gzCvlcIZVoM+14hlGcQ9r1Cbg2YqgJTvu7OBuAHhrnPFXts37rTIMVeBz0u9nponuF9O8LtLQU1YBD5uju7/NIdSfPYvnWnQYq9Dnpc7PXQPFefPxxubyko02LY9wqhPIOw7xVCmRbDvlcI5RmEfa8QyrQY9r1CKM8g7HuF3BowVQXmBmuvltnAfIeRW8TuSP59zWMkaBr/OblF9+3pgsZ13nkLuL2loAYMsvkmG2SWl+8w/jq47I7k39c8RoKm8Z+TW3Tfni5o3AF7d4bbWwrKtBj2vUIozyDse4VQpsWw7xVCeQZh3yuEMi2Gfa8QyjMI+14htwZMVYG59cbrZDZONjAru7GY/5w7jTveft4e57Mfu8/Z4xH/OfsWjdu77XZwe0tBDRhk1x23ziyzsMPYj23+c+407nj7eXucz37sPmePR/zn7Fs07siD9obbWwrKtBj2vUIozyDse4VQpsWw7xVCeQZh3yuEMi2Gfa8QyjMI+14htwZMVYE54sDsme6zG5pl30fj/PtB88hjNF2x5+xpNPfRc/5juWD/VcP6wO0tBTVgkGsuGGEtu7BD2dDzQfPIYzRdsefsaTT30XP+40YrLG+e/edVcHtLQZkWw75XCOUZhH2vEMq0GPa9QijPIOx7hVCmxbDvFUJ5BmHfK+TWgKkqMOWKAft13DGzkbKh+Q5j3+aDyEPT2c+749DzPvQact9WbDqfP26F5ZczIw/sDLdVAzVgELliwHGD98ssu7AD2bc+f5pi09nPu+PQ8z70GnLfVmw6nz9uxUYrmEkTRsJt1UCZFsO+VwjlGYR9rxDKtBj2vUIozyDse4VQpsWw7xVCeQZh3yvk1oCpKjB9FwztaVo0bWJWzFTSbgcqdeuzxxebxudOg+77j9GtO261lVc0XZtvbaac1BdunxZqQI0Hb77AdO/UwjRuvGJmnXAnLHbrs8cXm8bnToPu+4/RrTturTVWMwP362peemQK3D4tlGkp7HtZKE8N9r0slGkp7HtZKE8N9r0slGkp7HtZKE8N9r0stwZMZYHpu3/84eb6UQdmOs5WuTDy/MfurXvffhw0jT1Obovd96f15Z//kzlsz5bmplMHhD5Fggs1YDl+eOt+8+rU682A3l1r1xF1LvvWvW8/DprGHie3xe770/r85+UcYmeOPMy8/fRNoU+R4EKZarHv4Uy12PdwrhrsezhTLfY9nKsG+x7OVOuP3vfcGjDVBeYjFw4x+7TdrjaQbFhZ6L49zh2P7rvTuOMQNL3/eLlllzXD+3aC2xIGasBy/PrBI2bIoH28dfPZncy9b49zx6P77jTuOARN7z9efrnlzDXjw50eAUGZarHv4Uy12PdwrhrsezhTLfY9nKsG+x7OVOuP3vfcGjC1BaZ09B6tmnohZIMp5I9zb/37xcbbzxd7Do1zueP9eYRcbgttU7lQA2pJRz/0wB7W+gV3Onsaex53vP18sefQOJc73p9HyOW20DaVC2Wqwb7HvhcVylSDfY99LyqUqQb7HvteVG4NmNoC84DOO+VC8MOoez9onDte7vuP/fvuY3se9Jw9Hk3jP5avnscctDvcrnKgBtQaduQBufXBHdCGxrnj5b7/2L/vPrbnQc/Z49E0/uPlllvW3DhxDNyucqBMNdj32PfQdpUDZarBvse+h7arHChTDfY99j20XeVwa8BUFphy4frshvsB5G+LjXPH24pN4453x9mKvY7Lf51GKyxnrhy2H9w+LdSAGnLh+uz6FXYouS02zh1vKzaNO94dZyv2Oi7/dRqv1Mg8c9+VcPu0UKalsO9loTw12PeyUKalsO9loTw12PeyUKalsO9loTw12Pey3BowdQXmX0b3M40brZDZcD+8ure2YtOgaW2lppPxPnecO519a4/f6M+reztNo+3UQA1YyhtP/sWssnLjzDrkO5R7ays2DZrWVmo6Ge9zx7nT2bf2+C0328jbaRptpwbKNAj7Xh7KsxT2vTyUaRD2vTyUZynse3ko0yDse3koz1LY9/LcGjBVBaack0tOlZDd8Cz7vv3YvS1G81r2fbm177vP2/c10w3stivcVg3UgEHknFxyqoTsOhR2Jvexe1uM5rXs+3Jr33eft+9rpht9/EC4rRoo02LY9wqhPIOw7xVCmRbDvlcI5RmEfa8QyrQY9r1CKM8g7HuF3BowVQXmZcf3ym1sNjB033+Mbv376Hk0Tm7Rffux+7z72L+PphGNV1zB3HP2oXB7S0ENGOTJuy/LrUe2o6D7/mN0699Hz6Nxcovu24/d593H/n00jVh1lcbmi1fvgdtbCsq0GPa9QijPIOx7hVCmxbDvFUJ5BmHfK4QyLYZ9rxDKMwj7XiG3BkxVgdmr/Q6ZDfXDyt/aHajY83LfHm8/h6axx9mP/XHutJr50Hh5LPu3oO0tBTVgkKMP6ZVZZnAHKva83LfH28+haexx9mN/nDutZj40Xh7L/i1oe0tBmRbDvlcI5RmEfa8QyrQY9r1CKM8g7HuFUKbFsO8VQnkGYd8r5NaAqSowd9pig9zG+kGVJtPZ86D57fv246Bbnzy22ePs6f1x7mO532+3neH2loIaMEjH1v5RgMU7k0ums+dB89v37cdBtz55bLPH2dP749zHcv+ko/vB7S0FZVoM+14hlGcQ9r1CKNNi2PcKoTyDsO8VQpkWw75XCOUZhH2vkFsDpqrA7N1hB2/jshubZ4+zb9F0QdO4j232PPY4e7z7nH2L7vuPRw3YDW5vKagBgxx7WG9ruYWdxx9n36LpgqZxH9vseexx9nj3OfsW3fcfX3/JKLi9paBMi2HfK4TyDMK+VwhlWgz7XiGUZxD2vUIo02LY9wqhPIOw7xVya8BUFZj/PP9w07dzM9O0ybpm43XWMButs7pH7vuP7Vt3vH3fv22ybva+z3/OHWezx7vTFLvvarLummaHzdY3x/Rq553AFm1vKagBg3z/1j/N8CF9TYtmTc3Wm29sttpsI4/c9x/bt+54+75/u80WTbz7Pv85d5zNHu9OU+y+q+mWTUy7FjuYi8Yd453AFm1vKSjTYtj3CqE8g7DvFUKZFsO+VwjlGYR9rxDKtBj2vUIozyDse4XcGjBVBSYVQg1IeihT0kF5kh7KlHRQnqSHMiUdlCfpuTVgogUmWgHSQ/8BSAflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGLFlgtm/T0gw+ZJA5Y9xp5rxzzjJnnznODD/xeLNn991Ni112gvP4UAOSHmpA0kF5kh7KlHRQnqSHMiUdlCfpoUxJz60BAwvM3Tt3MOefe7a5bspkc/21UwpcfeUV5uCD+gcWmagBSQ81IOmgPEkPZUo6KE/SQ5mSDsqT9FCmpOfWgEULzFbNdzannTq6tqA89+yzzLFHDzUjh51oJl19lTdu8jVXmx7ddoPzC9SApIcakHRQnqSHMiUdlCfpoUxJB+VJeihT0nNrwKIF5r5772munTzJKyRPHX2KaduquTdevrE8aEA/M2XS1d7zUnS68/pQA5IeakDSQXmSHsqUdFCepIcyJR2UJ+mhTEnPrQGLFpijRo7wikv5tnKvHt1My12bmXatW3hat9gFzuNCDUh6qAFJB+VJeihT0kF5kh7KlHRQnqSHMiU9twaEBab8PH7G6WO9AnPC+PNM7332MuNOO9Xb71IKzgvOP9ccMfhQ07ZVizrz2lADkh5qQNJBeZIeypR0UJ6khzIlHZQn6aFMSc+tAWGBKUeOX3zhBK/AlKLy6isv9+5PmXRNwQE/8tN50LeZqAFJDzUg6aA8SQ9lSjooT9JDmZIOypP0UKak59aAsMDs1L6NufLyibWF5FVXTDSHDBpoeu7Z3fQ7oI+5cMJ4b/x11042hxw0oM78PtSApIcakHRQnqSHMiUdlCfpoUxJB+VJeihT0nNrQFhgdmjb2lx2ycXZInJK3SKy1z571R5JfsrJI4ueqgg1IOmhBiQdlCfpoUxJB+VJeihT0kF5kh7KlPTcGhAWmPKzt5xQXQpI+Vl87z27FzwvB/r4BaicJ7PYz+SoAUkPNSDpoDxJD2VKOihP0kOZkg7Kk/RQpqTn1oCwwBQnHn9s7c/ggwb2K3hu7z33qP0GczS/wUwMakDSQXmSHsqUdFCepIcyJR2UJ+mhTEnPrQGLFpjdd+9SW0RecfllZkC/A7xzYe7bc09z8YUXeOPFwQP7w/kFakDSQw1IOihP0kOZkg7Kk/RQpqSD8iQ9lCnpuTVg0QJTHHbwQd5P5H4xaZN9M8fyKPJEoQYkHZQn6aFMSQflSXooU9JBeZIeypT03BowsMCUn74PPKCPueD888w1V13pFZtye+nFF5ohRxxm2rTcFc7nQw1IeqgBSQflSXooU9JBeZIeypR0UJ6khzIlPbcGDCwwfXLi9T2772567b2Xd+3xUoWlDzUg6aEGJB2UJ+mhTEkH5Ul6KFPSQXmSHsqU9NwaUFVghoUakPRQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOypP0UKakg/IkPZQp6aA8SQ9lSnpuDZhogYlWgPTQfwDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQFZYKYYakDSQ5mSDsqT9FCmpIPyJD2UKemgPEnPrQEDC8zdOrU3A/r1Lap/3/1N6xa7wHkFakDSQw1IeihT0kF5kh7KlHRQnqSHMiUdlCfpuTVgYIE59IjB5vprpxR13ZTJplP7tnBegRqQ9FADkh7KlHRQnqSHMiUdlCfpoUxJB+VJem4NGFhgDh92vFdITr7manPRhAvquPCC802Hdq3hvAI1IOmhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGjCwwBw96iSvwDz/3LNN+7atTPs2LetosctOcF6BGpD0UAOSHsqUdFCepIcyJR2UJ+mhTEkH5Ul6bg1YtMCUwvG0U0d7BeYZ406D05SCGpD0UAOSHsqUdFCepIcyJR2UJ+mhTEkH5Ul6bg1YtMBs26q5982lFJhjR59iDh000JyZKTQvuehCc8bpY83AfgeYlrs2g/P6UAOSHmpA0kOZkg7Kk/RQpqSD8iQ9lCnpoDxJz60BixaYHdu1MZddcpFXYE6ZdI13Kwf1yK1/X35C51HkyUENSHooU9JBeZIeypR0UJ6khzIlHZQn6bk1YNECU05RdM1VV2YLzMnXmJHDT/ROTXTYIQeZSy/OFp7ioP4HwvkFakDSQw1IeihT0kF5kh7KlHRQnqSHMiUdlCfpuTVg0QJTDuoZfsLx5uQRw80hgwYW/By+z149zKSrs8XnqJNGFD3QBzUg6aEGJD2UKemgPEkPZUo6KE/SQ5mSDsqT9NwaMPAgnzatmnvcfS1bNd/ZXHLRBK/AlP00i/1MjhqQ9FADkh7KlHRQnqSHMiUdlCfpoUxJB+VJem4NWLTA7L57Z3PB+ed5BvQ7oOC53Tt3MFdePtErMMeOHsVvMBOCGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza8CiBWaXTu3N1Vde7hWR8m1lr3328grJzh3bmdGjTvbGiyFHDIbzC9SApIcakPRQpqSD8iQ9lCnpoDxJD2VKOihP0nNrwMCfyI8eekRtITnp6qvMpZdc5H1z6R9NPmH8eaZD21ZwfoEakPRQA5IeypR0UJ6khzIlHZQn6aFMSQflSXpuDVi0wBSyb+WRhx9mrr7yitpC0ycnYZcjzdF8PtSApIcakPRQpqSD8iQ9lCnpoDxJD2VKOihP0nNrwMAC0ycnXe+1915m0MB+pm+f3qZzh7ZwOhdqQNJDDUh6KFPSQXmSHsqUdFCepIcyJR2UJ+m5NaCqwAwLNSDpoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqQBWaKoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03Bow0QITrQDpof8ApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyJD2UKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPyrJZZnz1t5n3/lln46+dm0azvzeI5MzK335kFv3xq5n7zmpn1yRNwvmpCmZIOypP0UKakg/IkPZQp6bk1IAvMFEMNSDooz0qb/cXzXiFpapaaoKFm6SKz8LfPvUIUvU41oExJB+VJeihT0kF5kh7KlPTcGpAFZoqhBiQdlGflTDULfvkkUznW5EpI3SCFpnzTiV+zslCmpIPyJD2UKemgPEkPZUp6bg3IAjPFUAOSDsqzIqY9YRbP+TFXMoYbpDiFr11BKFPSQXmSHsqUdFCepIcyJT23BmSBmWKoAUkH5VkJi2Z9mysTow3zZ3wAX79SUKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOyjNp8394N1cexjDU1Jg5X74Al1MJKFPSQXmSHsqUdFCepIcyJT23BmSBmWKoAUkH5ZmkWZ88ZWqWLMxVh/EMS+b9CpdVCShT0kF5kh7KlHRQnqSHMiU9twZkgZliqAFJB+WZpPk/vp8rC+Md5nz5Ilxe0lCmpIPyJD2UKemgPEkPZUp6bg3IAjPFUAOSDsozSfJtYxLDwl+nw+UlDWVKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDwTM+3xkue6DDssmf8bXmbCUKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOyjMps6c/kysH4x9kv060zKShTEkH5Ul6KFPSQXmSHsqU9NwakAVmiqEGJB2UZ1Lkij1JDXLydbTMpKFMSQflSXooU9JBeZIeypT03BqQBWaKoQYkHZRnUmZP/3euHIx/qFm8AC4zaShT0kF5kh7KlHRQnqSHMiU9twZkgZliqAFJB+WZmGlTTc3SxbmSMN5hybxf8DIThjIlHZQn6aFMSQflSXooU9Jza0AWmCmGGpB0UJ5JWjxnRq4kjHdY8PM0uLykoUxJB+VJeihT0kF5kh7KlPTcGpAFZoqhBiQdlGeS5n33Zq4kjHOo8Q4gQstLGsqUdFCepIcyJR2UJ+mhTEnPrQFZYKYYakDSQXkmatpUs3Th7FxhGM8g1zWHy6oAlCnpoDxJD2VKOihP0kOZkp5bA7LATDHUgKSD8kza3K9fNnIN8TgGOT3R7M/+BZdTCShT0kF5kh7KlHRQnqSHMiU9twZkgZliqAFJB+VZCfNnfJArESMMNUszxeor8PUrBWVKOihP0kOZkg7Kk/RQpqTn1oAsMFMMNSDpoDwrZf6MD6VKzBaLZQ5yNPrcb16Dr1tJKFPSQXmSHsqUdFCepIcyJT23BmSBmWKoAUkH5VlJc7951TuHZTnDkgW/m9mfPwdfr9JQpqSD8iQ9lCnpoDxJD2VKem4NyAIzxVADkg7Ks9IWz/kxVzrqhgU/fQxfpxpQpqSD8iQ9lCnpoDxJD2VKem4NyAIzxVADkg7Ks9IWz/05VzrqhoW/fgZfpxpQpqSD8iQ9lCnpoDxJD2VKem4NyAIzxVADkg7KM2mzPnnCzP/xvUxh+ZNZunh++UeU1yw1SxfNNYtmfW/mffc/79RHaDmVgDIlHZQn6aFMSQflSXooU9Jza8CyCszdOncwe+7R1bNH191My12bwel8qAFJDzUg6aA8kzTnq5eyRWWMw5L5M73rnKPlJQ1lSjooT9JDmZIOypP0UKak59aA6gJzz+67mysvn2iuv3aK59rJk0yXju3htD7UgKSHGpB0UJ5JkavtJHUtcjl5+6xpT8DlJgllSjooT9JDmZIOypP0UKak59aAqgKzbavm5uwzx9UWlywwKwM1IOmgPJOy8LcvcuVgMsO879+Gy00SypR0UJ6khzIlHZQn6aFMSc+tAUsWmC122ckcefih5ropk82USdeYiy+cwAKzQlADkg7KMynlHsxT7rDgl0/hcpOEMiUdlCfpoUxJB+VJeihT0nNrwJIFZg/rp/FRI0eY4ScezwKzQlADkg7KMykLf52eKwWTGbwDfsByk4QyJR2UJ+mhTEkH5Ul6KFPSc2vAwAKzTctdzeljx3gF5aUXX2R269TenHDcMSwwKwQ1IOmgPJMi1wyXa4cnMciBPr9PexwuN0koU9JBeZIeypR0UJ6khzIlPbcGDCwwBw3o5xWS4qD+B3rjWGBWDmpA0kF5JmnOF/8xSxfOyZWF8QxyuqNZnz4Nl5c0lCnpoDxJD2VKOihP0kOZkp5bAxYtMDt3aGsuu+Rir5gce+po06r5zt54FpiVgxqQdFCeiZs21cz77k3vko9RBrkC0NyvX8HLqBCUKemgPEkPZUo6KE/SQ5mSnlsDwgJTDuzx97W86oqJZo+uXWqfY4FZOagBSQflWRlTIxeYi2Z+BV63slCmpIPyJD2UKemgPEkPZUp6bg0IC8zdO3fwCkgpJC+aMN4cPfSIWuedc7Y3Xo4qlyL0iMGH1n676UINSHqoAUkH5VkJc79+OVcmhh9qli6p2k/jPpQp6aA8SQ9lSjooT9JDmZKeWwPCArPbbp28IlLjiomXmXatW9R5DYEakPRQA5IOyrMSlsz7JVcmRhvkyHT0+pWCMiUdlCfpoUxJB+VJeihT0nNrQFhgdu7Qzjux+tlnnlGHFJR+cXn+uWeb0aNO8o42R6+DGpD0UAOSDsozaXI6odiGmqVm9ufPweVUgpsn6aE8SQ9lSjooT9JDmZKeWwMWPcinmJNGDPOKS+6DmTzUgKSD8kzSrM+eNjWLF+Sqw3iGJfN/9Q4cQstLGsqUdFCepIcyJR2UJ+mhTEnPrQHLLjBHDj+RBWaFoAYkHZRnYjJFoJxSKImhGlfxEShT0kF5kh7KlHRQnqSHMiU9twYsu8Ds2K6N6b57Z9Ntt86m5a7N4DQ+1ICkhxqQdFCeSUn2WuQ1vBZ5PYPyJD2UKemgPEkPZUp6bg1YdoFZDtSApIcakHRQnklY+MtnuUIwwaEmU2RW+HKRKFPSQXmSHsqUdFCepIcyJT23BmSBmWKoAUkH5RmvqWbhb5/nKsAKDFJkfv8WWI9koExJB+VJeihT0kF5kh7KlPTcGpAFZoqhBiQdlGdspk01i37/Olf5VXKoMfNnvI/XKWYoU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflGYtpj5tFs77PFXzVGRb8PA2vW4xQpqSD8iQ9lCnpoDxJD2VKem4NyAIzxVADkg7KMw7V+eay7jD/x/fg+sUFZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPKOa++3rufIuBUPNEjN7+r/hesYBZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPKNaPLu6P427w4KfPoLrGQeUKemgPEkPZUo6KE/SQ5mSnlsDssBMMdSApIPy1Jr9+bPeT9BylPiimV/VqlkS75V6og5LF84uWD+5frmcM3PWp0/D7SoHypR0UJ6khzIlHZQn6aFMSc+tAVlgphhqQNJBeZYy67N/mcWzf8iUbjXZCq6+DjVLvWLz92lPwO3UQJmSDsqT9FCmpIPyJD2UKem5NSALzBRDDUg6KM8gUlwuXTQvV6E1jGHJvF+8o97R9paCMiUdlCfpoUxJB+VJeihT0nNrQBaYKYYakHRQnkHkJ+aGOMz/4V24vaWgTEkH5Ul6KFPSQXmSHsqU9NwakAVmiqEGJB2UZ5Cli+bmSrKGNSya9R3c3lJQpqSD8iQ9lCnpoDxJD2VKem4NyAIzxVADkg7KM8iS+TNzJVnDGhbO/BJubykoU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflGWTeD+/kSrIGNNQsNXO+fAFubykoU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflWYqclqjBDJniUopmtJ0aKFPSQXmSHsqUdFCepIcyJT23BmSBmWKoAUkH5akx9+tXzOI5M0xNzZJcpVa/hpoli8yi378xs794Hm6fFsqUdFCepIcyJR2UJ+mhTEnPrQFZYKYYakDSQXmWY9a0J8zsz5/LFGvf5kq3NA81ZsFPH5vZ058JfVoiF8qUdFCepIcyJR2UJ+mhTEnPrQFZYKYYakDSQXmWZ6p3gEy9GWpqzPwIP4m7UKakg/IkPZQp6aA8SQ9lSnpuDcgCM8VQA5IOylNvqln0+9e5yq1+DXKJS7xN5UGZkg7Kk/RQpqSD8iQ9lCnpuTUgC8wUQw1IOihPLbnMYv0dasy8796E21UOlCnpoDxJD2VKOihP0kOZkp5bA7LATDHUgKSD8tSY9/3buUKtHg81S0KfnsiHMiUdlCfpoUxJB+VJeihT0nNrQBaYKYYakHRQnqXM/vxZU7O0fh497g5yZSI5UAltpwbKlHRQnqSHMiUdlCfpoUxJz60BWWCmGGpA0kF5liKnJ2pIw4JfPoHbqYEyJR2UJ+mhTEkH5Ul6KFPSc2tAFpgphhqQdFCeQeZ89VKuLGs4Q83SxWbWp0/B7S0FZUo6KE/SQ5mSDsqT9FCmpOfWgCwwUww1IOmgPIMs/O2LXFnWsAbZpxRtbykoU9JBeZIeypR0UJ6khzIlPbcGZIGZYqgBSQflGWTx3J9zJVnDGhb88inc3lJQpqSD8iQ9lCnpoDxJD2VKem4NyAIzxVADkg7KM8iCX6ebmpoaT0Ma5n3/FtzeUlCmpIPyJD2UKemgPEkPZUp6bg3IAjPFUAOSDsozyKxPnjALfvnMLJk/0yxZMNssXTinHpttlsz71cyf8UFm26bW2VYNlCnpoDxJD2VKOihP0kOZkp5bA7LATDHUgKSD8iQ9lCnpoDxJD2VKOihP0kOZkp5bAyZaYKIVID30H4D0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0AWmCmGGpD0UKakg/IkPZQp6aA8SQ9lSjooT9Jza0BVgblbp/am1z57mf1772v223dv0333zqbFLjvBaW2oAUkPNSDpoUxJB+VJeihT0kF5kh7KlHRQnqTn1oCBBWbb1i3M8cceba6YeJm5dvIkc/21U8x1Uyabq6+83Jxy8kjTsV1rOJ8PNSDpoQYkPZQp6aA8SQ9lSjooT9JDmZIOypP03BqwaIHZqvnOZtRJw72iUkyZfI258vKJtYWmGHfaqaZ1i13g/AI1IOmhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGrBogblH1y61xeQ5Z55hOnds5xWTXbt0MhdNuMAbf921k83unTvC+QVqQNJDDUh6KFPSQXmSHsqUdFCepIcyJR2UJ+m5NWDRAnNgv77m8ssuNRMvvcTsvdceBc8ddsig2m8xZZ9M+zkbakDSQw1IeihT0kF5kh7KlHRQnqSHMiUdlCfpuTWg6iAfW9tWzb2fxqW4nHT1VaZzh7ZwOoEakPRQA5IeypR0UJ6khzIlHZQn6aFMSQflSXpuDagqMOXn8mEnHGdGDj/RnH/u2bkDfa4wRww+NPBoctSApIcakPRQpqSD8iQ9lCnpoDxJD2VKOihP0nNrQFWBeVD/A2t/EvedPnaM6dql+P6XAjUg6aEGJD2UKemgPEkPZUo6KE/SQ5mSDsqT9NwaUFVg7tl9dzPixOPNSSOGmTPHnWamTLrGKzInXnqx6d61C5xHoAYkPdSApIcyJR2UJ+mhTEkH5Ul6KFPSQXmSnlsDlr0Pppy+aPChB9ceYS4/mxf7mRw1IOmhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGrBogdl3/97m6CFHmiMOO8S0a9Oy4Dm5ks9VV1zuFZjnn3tO0XNhogYkPdSApIcyJR2UJ+mhTEkH5Ul6KFPSQXmSnlsDFi0wjz/uaK+AlAN6DjvkoNpvKeX28EzRed2U7DeYp4891ftW051foAYkPdSApIcyJR2UJ+mhTEkH5Ul6KFPSQXmSnlsDFi0wZb9LOVLcLzLPOuN0c+Lxx2Zux3mPZbz8TN7vgD5wfoEakPRQA5IeypR0UJ6khzIlHZQn6aFMSQflSXpuDRi4D2a/vn28E61LMem68vLLvH0xW+7aDM4rUAOSHmpA0kOZkg7Kk/RQpqSD8iQ9lCnpoDxJz60BSx7kIydSP/Tgg8zJI4ebM04/zZxy0ohMYTnI7NapPZzehhqQ9FADkh7KlHRQnqSHMiUdlCfpoUxJB+VJem4NWLLAjAI1IOmhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGpAFZoqhBiQ9lCnpoDxJD2VKOihP0kOZkg7Kk/TcGjDRAhOtAOmh/wCkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwOywEwx1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwP+YQrMWZ89beZ9/5ZZ+OvnZtGs783iOTMyt9+ZBb98auZ+85qZ9ckTcL5qQg1YLU9PGmXeeuSv5vPX/s98/9HrZsb098x3H75qPv3vVPPafdeYJ644Ac5XLShP0kOZVgv7Xnh834uGfS889r1o6lvfE24N2OALzNlfPO91alOz1AQNNUsXmYW/fe79p0CvUw2oASvt+ZvOyXTq18zSJYtzSeFh0YK55vPXn/b+U6DXqTSUJ+mhTCuNfS88vu9Fw74XHvteNPW17wm3BmzABebUzF9Kn2R6cU2uOXSDdHr5qwu/ZmWhBqyUqZccbT556dFMHkv8ZHK3Msh9V3aQTv/WIzfC16wklCfpoUwrhX0vCr7vRcG+FwX7XhT1ve8JtwZsmAXmtCfM4jk/5uIPN8h/FPjaFYQasBKemHi8+fGTt3JJyJDvzMH3/cc13n+Uxy4+qs5rVwrKk/RQppXAvhcB3/ciYd+LgH0vkobQ94RbAzbIAnPRrG9zoUcb5s/4AL5+paAGrIRvP3gll4AM+Q5ceN8f/PH2uOzwwdP3wNevBJQn6aFMK4F9Lzy+70XDvhce+140DaHvCbcGbHAF5vwf3s1FHcNQU2PmfPkCXE4loAZM2rtP3J7beBnczu127GK3MtR4X/W/cOt4uJykoTxJD2WaNPa98Pi+Fw37Xnjse9E0lL4n3BqwQRWYsz55ytQsWZgLO55hybxf4bIqATVgkp66crhZOHdWbsvtTi2DfV8G//ng6X79+hO4rKShPEkPZZok9r3w+L4XDfteeOx70TSkvifcGrBBFZjzf3w/F3G8w5wvX4TLSxpqwCS9/39/y22xDHYnLuzA2cHt4Pa09n1jXrx9AlxeklCepIcyTRL7Xnh834uGfS889r1oGlLfE24N2KAKTPnLJ4lh4a/T4fKShhowSfKXT76jylCsA7vT2M/5t/n70199Ci4vSShP0kOZJol9Lzy+70XDvhce+140DanvCbcGbDgF5rTHM7kGn3cr7LBk/m94mQlDDZiUxyceZ5YuXpTZWtRx7cHvyPbz7mN/yN7/7bvpcJlJQnmSHso0Kex7EfB9LxL2vQjY9yJpaH1PuDVggykwZ09/xgs2iUH2MUHLTBpqwKQ8c8Pp/tYWIUOx+zKg57JkHxO0zCShPEkPZZoU9r3w+L4XDfteeOx70TS0vifcGrDhFJhfPC8pJzLIiWDRMpOGGjApz990dm5rZbA7rT/4nVcG+9YdX5ecCBYtM0koT9JDmSaFfS88vu9Fw74XHvteNA2t7wm3BmxA32D+OxNsMkPN4gVwmUlDDZiUf197qr+1Fn+w78vgP7Zv3XH5YcGcmXCZSUJ5kh7KNCnse+HxfS8a9r3w2PeiaWh9T7g1YAPaB3Nq5q+e4Gt3hh2WzPsFLzNhqAGTMvXSo83iBfMyW2t3Vr8Tux0ZTWMP9rga88tXH8FlJgnlSXoo06Sw70XA971I2PciYN+LpKH1PeHWgA2nwMxYPGdGLuB4hwU/T4PLSxpqwCTN+Oyd3BbnO2rd+/5jGdBzLmOm/edBuLwkoTxJD2WaJPa98Pi+Fw37Xnjse9E0pL4n3BqwQRWY87570ws33qHG25kZLS9pqAGT9ObDN3jb63bW/K072NP4g/24xtTULDXPXH8aXF6SUJ6khzJNEvteeHzfi4Z9Lzz2vWgaUt8Tbg3YoApM+cp+6cLZuaDjGeQaq3BZFYAaMElTLz3GzP75u9yW+x3Z7dBBj93xxnz7/itwWUlDeZIeyjRJ7HsR8H0vEva9CNj3ImlIfU+4NWDDKjAz5n79ciZnO/Twg5wqYfZn/4LLqQTUgEl7+W+Xmpql9rnN7I6M7suAnsueKuFfU0bD5SQN5Ul6KNOkse+Fx/e9aNj3wmPfi6ah9D3h1oANrsAU82d84MUeaahZmvmP8wp8/UpBDVgJH/z7XgkgRwb/VgZ3nH2bt3TJYvPKPZfD168ElCfpoUwrgX0vPL7vRcO+Fx77XjQNoe8JtwZskAWmmD/jw1zw5Q9yZNzcb16Dr1tJqAEr5cNn/pH5o9TuwP5gj7PJkL1dvHC+ee0fV8PXrRSUJ+mhTCuFfS88vu9Fw74XHvteNPW97wm3BmywBaaY+82r3vm0yhmWLPjdzP78Ofh6lYYasJJevfcK73xahR3aHuxx2fu///iVee6vZ8LXqySUJ+mhTCuJfS88vu9Fw74XHvteNPW57wm3BmzQBaZYPOdHrxG0w4KfPoavUw2oASvtx0/fziXjd3i/g9u3+fsfP3c/fJ1KQ3mSHsq00tj3wuP7XjTse+Gx70VTX/uecGtAVYHZqvnOpnOHtma3zh3Mbp3am47tWpsWu+wEp7WhBqy0xXN/zjWEblj462fwdaoBNWCl/fyF+7NHYefO32bvf/bKE/B1Kg3lSXoo00pj3wuP73vRsO+Fx74XTX3te8KtAQMLTCkie/bobk47dbS5+srLzXVTJptrJ08yl192iTn+2KO9QhPN50MNmLRZnzxh5v/4XqaT/2SWLp6faQO/QZRDzVKzdNFcs2jW92bed//zTsOAllMJqAGT9sQVJ5j3nrrT/DT9PTN/1q+ZOPyj2/wO7eeJb2VH47kzfzLff/S6+d+D13lXK0DLSRrKk/RQpklj3wuP73vRsO+Fx74XTUPpe8KtAQMLzF5772WuyhSW1187xSsuJ19zlVdgymMx7rRTTZuWu8J5BWrAJM356qVsB49xWDJ/pnfNVbS8pKEGTNJLd1xo5v/+S27L/QF1ajTOv7WfN2bmd59711xFy0sSypP0UKZJYt8Lj+970bDvhce+F01D6nvCrQGLFphSOJ595hleITnp6qvM4EMGme67d84UnXuaCePPry0y++7fG84vUAMmRc78n9R1UeVEsrOmPQGXmyTUgEmRM/9nr4sqg91p7c7r39pDsefy42f/9K154vLj4XKTgvIkPZRpUtj3wuP7XjTse+Gx70XT0PqecGvAogWm7G8phaUUkaeeMqpgn8v+fff3vtGU54475qiC+WyoAZOy8LcvcuEmM8z7/m243CShBkzKF2/8O7el0kl9/mA/dp/X3b796E1wuUlBeZIeyjQp7Hvh8X0vGva98Nj3omlofU+4NWDgN5j9DuhjBvbr631zaT/Xr2+f2gLz6CFHFDxnQw2YlHJ3LC53WPDLp3C5SUINmJSfv5AT5bodVQa5b493yYDGC3+oMZ/+t7Lbg/IkPZRpUtj3wuP7XjTse+Gx70XT0PqecGvAwH0wkfZtWprx557jFZdTJl2TKT67wOkEasCkLPx1ei7YZAZv52Ow3CShBkzK9FefzG0p6rDuYxnc52Tw79d97n8PXQ+XmxSUJ+mhTJPCvhce3/eiYd8Lj30vmobW94RbA5ZVYLZt1dycOnqUV1zKN5jHHDUk8HRFqAGTItcvleuYJjHITse/T3scLjdJqAGTItcvleuYFnZUe3A7sDudfyuD/bwxM7//3Dx+2bFwuUlBeZIeyjQp7Hvh8X0vGva98Nj3omlofU+4NaC6wGzXuoUZc8pJtcXlKSePNK1b7AKn9aEGTNKcL/5jli6ck4s4nkFOvTDr06fh8pKGGjBJ/7n5XDPnl+8zW213YLvj2o+LjfeH7P2fPn/fPD3pZLi8JKE8SQ9lmiT2vfD4vhcN+1547HvRNKS+J9waUFVgtm/byowdfUptcTl61Enet5loWhtqwMRNm2rmffemd/mpKINcjeCPeOF9OYfWmw//xbv8VHZwO7Lboe3HMmTHydUIshfeP6rOMioB5Ul6KNOkse9FwPe9SNj3ImDfi6Sh9D3h1oAlC8wOmeLy9LFjaovLk0cMM20UxaVADVgZUyN39kUzvwKvW1moASth6iVHmd9/+DKTgtuR3cHu7PZtjfnqrefha1cKypP0UKaVwL4XBd/3omDfi4J9L4qG0PeEWwMGFphypZ4zxo2tLS6HnXBc4InVXagBK2Hu1y9nc48w1CxdUrWv6X2oASvh5bsv81NwyIDu24+zw5JFC6r2Nb1AeZIeyrQS2PfC4/teNOx74bHvRdMQ+p5wa8CiBab8BH7muNO84lLIEePjzzvXnHv2mQXkPJgtd20GXwM1YCUsmeeeGT/cIEfJodevFNSAlfDLVx/nEpABd+bC+zLY02Tvy1Fy6PUrAeVJeijTSmDfC4/ve9Gw74XHvhdNQ+h7wq0BixaYu3Vqb66+6oraArMYKUJbNd8ZvgZqwKTJqQ1iG2qWmtmfPweXUwlu41WCnNogt/G5W3/Id+K69/3bwvFLFy8yz/31DLicpKE8SQ9lmjT2vfD4vhcN+1547HvRNJS+J9waMOAbzBbmiMMOMUOPPDyQXNWn2KmKUAMmadZnT5uaxQtyYcczLJn/q7cTM1pe0lADJunpSaPMgjkzc1sug92BbTLY9+2hcLpfv/m0KhffR3mSHso0Sex74fF9Lxr2vfDY96JpSH1PuDVgyYN8okANmJhMh5TTGyQxVOOKAgI1YFKkQ/40/b3cFtsdNt9xs4P92H7eHucP2fuf/ncqXGaSUJ6khzJNCvteBHzfi4R9LwL2vUgaWt8Tbg3YYArMZK+LWtPAr4t6lPK6qP4497EM7n3/cY2pqakxbz92M1huclCepIcyTQb7XhR834uCfS8K9r0oGl7fE24N2CAKzIW/fJYLNsEh02CVvnQVasD4HWU+e/nx3Eb6A+rEfgd2n0Pj/Nv8fTlC8H8PXgeWnwyUJ+mhTOPHvhcF3/eiYN+Lgn0viobZ94RbA9bzAnNq5q+oz3OBVmCQDv/9W2A9koEaME5y7q3PX3/a37iAW58M2vv+kB9fs3SpeevRm+C6xA3lSXoo0zix70XB970o2PeiYN+LoiH3PeHWgPW3wJw21Sz6/WsvxMoONWb+jPfxOsUMNWBcZP+Pr999sXab8rdB9+3H9uBOJ4N/336c+TfzhvH+03fDdYoTypP0UKZxYd+LgO97kbDvRcC+F0lD73vCrQHrZ4E57XGzaJZcv7N6w4Kfp+F1ixFqwDjIRfC//+j13Ja4nVMGzbhi42Xwb2Xwx9vPGzPtPw/BdYsLypP0UKZxYN+LgO97kbDvRcC+F8kfoe8JtwaslwVmdf6KqjvM//E9uH5xQQ0Y3VHgrygZ/Pv2rWacDOh5GfzH9vP+bY1576k7wfrFA+VJeijT6Nj3ouD7XhTse1Gw70Xxx+h7wq0B612BOfdb/6+AFAw1S8zs6f+G6xkH1IBRvX7fJFnx7PqXdRtEBvdWBnucTYYas2TxQvPv68bC9YwK5Ul6KNOo2PfC4/teNOx74bHvRfNH6XvCrQHrXYG5eHZ1v6Z3hwU/fQTXMw6oAaP6/uM3cmvudzoZCjthfvDH28/L4I73n7Nv0Th/yD//0bP/hOsZFcqT9FCmUbHvhcf3vWjY98Jj34vmj9L3hFsDprbAnP35s97X4XLE2qKZX9WqWRLvVQOiDksXzi5YP7mWqpy/K46L9qMG1Hr2L2d4X4fLEWtfvfV8rQVzfs+sNep4/jj7ORmCpvUH/7F9a0/n3vpDjZn983cF6zf9lSe983dFvWg/ypP0UKZa7Hs4Uw2+77Hvoe3SQnlqse+x76HtKodbA6auwJz12b8yfzH94AVRr4eapdkL9097Am6nBmrAUv41+RTzw7T/eUeOFR/kOZs/oPHocdBgTysDuu9PYz9XOMg1Vae/9pR5YuLxcDtLQXmSHsq0FPa9LJRnKXzfy0OZlsK+l4XyLIV9Lw9lWgr7Xp5bA6aqwJSOvnTRvNzmNoxhybxfvCPw0PaWghowiHT0eb//nFuy3aGCyBB03x/88UHj0HMyoGnc51zZ4ZevPvKOwEPbGwTlSXoo0yDse3kozyB83yuEMg3CvpeH8gzCvlcIZRqEfa+QWwOmqsCUr7sb4jD/h3fh9paCGjCIfN2dHfzO4nYgnwyax/atDPY0iAzaxzLYzxUbb8y7T9wGtzcIypP0UKZB2PfyUJ5B+L5XCGUahH0vD+UZhH2vEMo0CPteIbcGTFWBuXTRXG/jGtqwaNZ3cHtLQQ0YZO5vMzJLsztMsSHfkfL3NY8RGdB4IYN/K4N7355OBjzuuw9fhdsbBOVJeijTIOx7eSjPIHzfK4QyDcK+l4fyDMK+VwhlGoR9r5BbA6aqwFwyf2ZuAxvWsHDml3B7S0ENGGTm919kluZ2GPuxTQb7tth4/9Yd5w/2Y/c5f/Dnd8ng3spQOO7LN5+F2xsE5Ul6KNMg7Ht5KM8gfN8rhDINwr6Xh/IMwr5XCGUahH2vkFsDpqrAnPfDO97GNaihZqmZ8+ULcHtLQQ0Y5J3Hb80tVAbpKHanscng3vdv3fv+Yxm0z/m32vvoORlqzNIli80Lt46H2xsE5Ul6KNMg7Ht5KM8gfN8rhDINwr6Xh/IMwr5XCGUahH2vkFsDpqrAFBW9kH7SQ6ajy39gtJ0aqAGD+RfSdzuQfesP/jTFprOfd8fJYD9nk8G+9e/bQ7HpfDJkO/o7U28F21kaypP0UKbB2Pd8KM9S+L6XhzINxr7nQ3mWwr6XhzINxr5nc2vA1BWYYu7Xr5jFc2aYmpoluQ2vX0PNkkVm0e/fmNlfPA+3Tws1oMYr91xuZkx/zyxZtFDWJkcGza1PBv9WBjSNzx+C7vuP0W3huEXz55hv3vuvef6mc+D2aaA8SQ9lqsG+F77v8X0vC2Wqwb7Hvse+5w/2dOi2cFwcfU+4NWAqC0zfrGlPmNmfP5fpON96IaR7qDELfvrYzJ7+TOhTJLhQA5bjicuPN8/99Uzz7fv/rV1H1LkKb9379mP/1r3vjvMHdN+f1pcd5BxiHz//gHnm+tNCnyLBhvIkPZRpOdj3wuP7Hs5Vi30vPPY9nKvWH7nvCbcGTHWB+fvHU72ddevNkGmw+RG+nnehBizH1EuONl/+75ncyvmD3cnc+/4tGi+De9+dxh2HyGDf5sfXLF1q3nk83OkRXChP0kOZloN9Lwq+70XBvhcF+14Uf+S+J9waMMUF5tTMX1FfeyHUt0Eut4W3qTyoAbWko3/9zgu5NZLB7ljZzoVv/fsyoPH28zKg59A4d3DH+/PUeJfbQttUDpQn6aFMtdj3cKY6fN9DmWqx7+FMddj3UKZaf/S+J9waMLUFplzyqf4ONWbed2/C7SoHakCt6a8+Wbsu+Vv3ftA4d7w/2PdlQM+5tzLIfXs8mkaGmswfpUvNmw//BW6XFsqT9FCmWux7OFMNvu+x76Ht0kJ5arHvse+h7SqHWwOmssCUC9fX+6FmSehTJfhQA2rIhetzKwFui41zx9tDsWnc8TLY42wyBD22xxuzZPFC88Jt4U6VIFCepIcy1WDfC9/3+L6XhTLVYN9j32Pfs8kQ9NgeH73vCbcGTF2BOfvzZ03N0vp5JJs7yFUSZKdptJ0aqAFLefYv48yShQsyS/c7Drq1yRB0W4wM9q3LHtxx7nT2bX783F9/9HaaRttZCsqT9FCmpbDvZaE8S+H7Xh7KtBT2vSyUZynse3ko01LY9/LcGjB1BaacKqEhDQt++QRupwZqwGBHeadKyA75TuN2InxbjAzofrHn/KHY8/Z997bu/U9eehRsZ2koT9JDmQZj3/OhPEvh+14eyjQY+54P5VkK+14eyjQY+57NrQFTVWDO+eolbwMb0lCzdLGZ9elTcHtLQQ0Y5KU7L/KXmruVwb3vP0a3/n0Z3OdlcMfJLbovg//Yfd59LIM7zn9szOKF881TV42A2xsE5Ul6KNMg7Ht5KM8gfN8rhDINwr6Xh/IMwr5XCGUahH2vkFsDpqrAXPibXNez4Q2yfwva3lJQAwb54o1/Z5ZWqgMVe94f3Ps2f3DH2Y/9cf5gj3OnsR8XG2+8/VvQ9gZBeZIeyjQI+14eyjMI3/cKoUyDsO/loTyDsO8VQpkGYd8r5NaAqSowF8/92du4hjYs+OVTuL2loAYM8vOXH+WWiDpNMf6A7tvT+Pftx0G3/iCPbTK49/1bd3z2/qf/nQq3NwjKk/RQpkHY9/JQnkH4vlcIZRqEfS8P5RmEfa8QyjQI+14htwZMVYG54NfpRs4uLxrSMO/7t+D2loIaMMj01/7Pys/mD/59d5w9XdA0/uA/tslg3/r3ZXDv29P5t+i+DDXmrUdvgtsbBOVJeijTIOx7eSjPIHzfK4QyDcK+l4fyDMK+VwhlGoR9r5BbA6aqwJz1yROZvzw+M0vmzzRLFsw2SxfOqcdmmyXzfjXzZ3yQ2bapdbZVAzVgkCcuP8F89vITZuZ3n5vZP39v5vz6Q9YvOf59e5z7uM401uvYz7njbPZ4d5pi9x2y/r9+/Yn54Ol7vBPYou0NgvIkPZRpEPa9PJRnEL7vFUKZBmHfy0N5BmHfK4QyDcK+V8itAVNVYFIh1ICkg/IkPZQp6aA8SQ9lSjooT9JDmZKeWwMmWmCiFSA99B+A9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2tAFpgphhqQ9FCmpIPyJD2UKemgPEkPZUo6KE/Sc2vAelNg3nb6QebSY/c1E47a21wwtKd3Ky46eh9v/NXD+5h/nDcYzvv3cw4zl5/Q21x4dHYee34Zd/Exmdc4rpeZNGJ/c1+x1zj3MDPx+F618/uv4c2bWf6Vw/Yzt542EM4bFmrAuPzywcPm/+653Pz03kPwedfMjx41V503zFxzwQj4fBqhTEkH5ZkecpWOcFfqqBSUaRo8elEWei4tUJ6khzKNw8MXHul9jj404Uj4vEv62bADOpoRB3aCz6cRyjOsD5+7zTx+16XmoVsmmAdvvsC7ffjWCebR2y/yxj93/9Xmmzf+Aef96rW/e5/Pj9x2YZ35Zdxjd1xsnvjbpeaFByeZb/93H3yNr1//u3nqnonePDK/kPsyryz/mfuuNO8/cyucNyy3BqwXBeZdZx5sGq2wnFlmmWUCrbHKSub+8YcXzCudfIsN14bTI6tnXkOKyTCvseyyfzKTRx5QMG8UqAHjcsW5J3jrvOO2W3gdGU1ju/iMY8yf/vSnTDssb15/4gY4TdqgTKvp3nMONUP2aWPa7rCpabVtEzOw266x/1ESF5Rntc3/4R2zZMHv3rVyhdyXcWjaakOZVtvt4waZ9ddezSP30TRpgPKsti9fu9ecP2aI2adbW9OjSysz+viBsX84xwVlGocT9u/gfWbIZ6EUmmga2zG922U+M5Yxyy+3rLnhlH5wmrRBeYbxyYt3mcYrNSqoD5B11l7D/PDW/QXzypc58rmMpkf+vNbqXjHpvsZO25V+jeUybfPSw5ML5o3CrQHrRYF52fG9YDjILWMLP7ClWJTCCE1bzF9GF/5n+Of5h6tf4+zBPQrmjQI1YFzOPeWI2nVefrnlzDGH9q7TSX03XzHW64j+9IcP6AmnSxuUabVIH15rtca1GfpWarS8GXPQ7nCeakJ5xmX29GfMvG/fMHO/ec3M+uxpOI1r0e/fZIpKPMhzaB6XLEuWKcuWdUDTxAVlWm2nH9Kttt/JfTRNGqA8q+nJuy8z66+zVsH/W7Fy45XMjRPHwHmqCWUahyN6tqrd9uWWXdb07rBDnS9jfGMHdfW+cPGn79lmWzhd2qA8w5A+4297Ke89c0vBvPI5bGen8caTfyl4je/f+qf6Ne6+7uyCeaNwa8B6UWCOH7JXbRhjxowxkydPLnDkkUfWPv/XMf0L5v3bWYfUPjdw4MA68/qOPvro2umuG3VgwWvIfyL/uQMOOKDOvBMmTKh9Ps43btSAcblo3DG16+xrstG65m/XnuX99eNPJ1+pr7Ri9i+xddZZx7tdZeXGZvrLdxe8XhqhTKvhjnGDzKqNV/SyW3755U2vXr3MoEGDzCqrrJIdlynerxrWB85bLSjPqKSoWzz351xZmBtqasyimV+bWZ88AecR875/Kzdx8UGmQfMKeW1ZhizLHmRdkio0UabVxgKzfB/95w6z5uqrFv2/u0Jm3LP/vArOWy0o0zgc06tdbf/xrbvmquaswXsU7HYhu441Wj77i6P/mdG40Qrm7sxnsf16aYTyDOP+m8bXZlSqZnnzqb8WzPvZf/9W+5y2ZnnlsesKXkOKVP+5UjXLbVefXjBvFG4NWC8KzHOP2LM2jFdeeSX38ZAf/va3fINce3Lfgnnl53X/uSlTpuTmqDvcd999tdNdM2L/gteQfTj956688srcHPnhm2++qX0+zm+jUAPG5fpLRnnrK28Aw4YNMyussIL3WL6p3b9nJ/Ph87eb/zxwjVl9tewb6VZbbWU+++wzs8EGG3iP5eci9LppgjKthkHdm9dm++ijj+Z6jTHvvvuuWW211bznOjXbAs5bLSjPKGZ99i9Ts3hBbsvrDkvm/WJ+n4b3q5TnSg3e/GBeec2g+WWdtN+ilgNlWmnXZ/5Q3q/jjmbvttt5mm+zsdfXhNz3x8s0Mi16jWpAeVbL2BMHlfy/K++XaN5qQZnGYdSA3bztrfuZkX3/kt0u5LNzldxPw+5nhuwehF43TVCeYfz9hnO9bRalapaXH722YN5PX7qr9jltzSKf1fZryD6c/nOlapY4v4V3a8B6UWCec3iP2jBQY9199921z2+50Z/N9putX6tpk3Vrn7v22mtzc9Qd/vnPf9ZOJ/uY2K+x7Sb515Dq3x3sxho9cDe4DWGgBozLvdef463vGmusYRYtWmReffVV06JFi9rtWGuN1cx666zp3V933XXNBx984G3ruHHjvHFbbLqhd6AQeu20QJlWQ4edNvcy22677bwM7aF///7ec7JfHJq3WlCeUXjfIJYYiu1PWbNkYW6K4oNMg+aV1yw1yLqheaNAmVZai6ZNvL6lIdOi16gGlGe19N4zu99h0P/dzZqsD+etFpRpHPzP4WKfGautvKJZc9XsbkDoM2PDP6/uHSiEXjstUJ5h+J+volTN0mz7LU3b5tvXatGsae1z2ppF9tm0X6PVLtvWPleqZvnLZaPhNoTh1oD1osCU/Rr9MFBjPfnkk7XPB7nxxhtzc9QdnnnmGTiPC72G3Vij+neB2xAGasC4yFFksr7yV+j8+fO97ViwYIE55ZRTardFyE9BL7zwgve8DJ9//nntX67ynwi9dlqgTKuhR6vsG8aaa65pZs6cmUvSmCVLlphdd93Ve26rzB9GaN5qQXlGUbNkUW6riw+L58yA8y5dODs3RfFBpkHzymuWGmTd0LxRoEwr7cQDOnrfJq24wvKeFXI/Wwq574+XaWRa9BrVgPKslkMPzH72BP3f3XmHreC81YIyjYOcLcXrOxE+M6RIRa+dFijPMGS/Rj+PtNcs1108Cm5DGG4N2CAKzNmzZ5sePXqYzTbbzGy44YbeV/Jy26RJE2/clltuaXbeeWcv1GLD3LlzTc+ePc3mm28OX2ObbbYx3bt3N1988UVujvxgN9ZJ/TrDbQgDNWBcXnv8Bm99l112WfPjjz+ab7/91owdO9astVZ+Z3Z5U7j//vtzW5kfZJ8Oeb5N8+3M6cMPMccP7mNOOLyPOfWEQd6pjOQ0CMVOnVBJKNNqsL+B79Kli3n++efNW2+9ZQ466KDa8Ufu3RrOWy0oT9esT//PzPnyBdV+jJphyfyZcN6Fv07PTVF8kGnQvPKamgHNa5NtlG2VbUbPu1Cm1fDoRUPMIxdmjT24a21/k/v+eJkGzVstKM9qsb+JKvZ/97zRR8J5qwVlGocbTjnQ294onxnbbbqeOWSPFqZPxx1Nn047ersPyamMLj5m36KnCKwklGcYpQrMNNUsUy48CW5DGG4NWD8KzBI/kftDTU0NVM6A5hdBg91YI+tJgSmnUZD9isSBBx5Yu9O6aNSokbdz8RtvvJHbwsLhxRdf9Obzp0dWXaWx6dm1jbnjmnFmxrsPwnVIGsq0GmQH+D1b53/2cDXbcgPz4AVHwHmrBeXpm/35c7lvBvP/L5YunGPmffc/OL1Yujj7jUfQsGjWd3BeKeqWLpqXm6ruIM8VK/zkNUsNsm5oXiHbJNuWH2q8bZcM0PQ+lGm18SCf8skBj4P75Y8BcHVq06xq72/FoEzjIMczyP6WSX1mNF5xBdNm+03NuEO7V+39EOUZxj0lCkx/QLWGKGdA84ugwa5ZJl84Em5DGG4N2CAO8qn2UFBgHlg/Cszv3ryvznm6Vl55ZXPccceZadOm5bYMD9J5BwwYYPbYYw/vSDY5Sk72s5G/ZuVxt27dCv6q3XTj9b1O/PP7upO6xwVlWi3yTZH89W7nLdZebeWip/qoJpSnmP3F84E/d8+f8QGcb8Evn+amKD7IKYTQvGL29H+bJfN+zU2ZH2ScPIfmEfKapQZZNzSvbEuxYenihV4WaD6BMq02Fpjh/PrBI96vNfb/W7HBumsXPbVbNaFM43Df+YPrnI86qc+M9dda1fuyRntS97igPMModZBPtQe7Zpk04Q9eYI4f2rM2jFtvvdW89tprqfLYY4/Vrl99+Yl86p2X1J4na+211/b+o8tPHnENso/O448/7v2l6+9/Izsv/9c5Yi5JKNNqkBOs77bLVrV9ZPXVV/d+xvAf77jFBubmUwfAeasF5SlQkVcwZD5IUMEnpwoK+rl64cwv68yD2Kc5kvtoGpe8drFB1mnWtLqnSJJtkG0pNsgH5uK5RY5cz0CZVhsLzPLJCdb79coePS3c/7sdWu1o3vnXzXDeakGZxuGSY/et/RayUp8ZcpCue2aYJKE8w3jAOk1R2muWP/xP5LJ/hh9G2p0yIP1Hkcsbovz1LevbsmVL88svpU8DE2WQU3rIviKyvMaNVzQ3XX4qXK+4oUwr7fwhe5l118j/lCRHXX788cfmp59+Mr17964dLwdaDO/bqeB8ctWE8pT9EDXD/J8+hPNLIbfw18/qfAMq49D0SM2S/KmO5D6aBpFl2IOsg4xDxaWQbdAMxfY/RZlW05ST+prOO+ev7CH3ZRyattpQntXwzxvPNxtvmD+DSLH/u3Iqt2vGDy84f3A1oUyjkj+A5dcW2d5Kf2bIgWinDqrMxShQnmHIcQh+/0i7Gy49BW5DGG4NWC8KTPkLptT+G2khJ5lF2xAGasCo5PxYOzbNnjZHzuMm/5ErMSxdutRcf/31mQKzsXdVoKvPHw7XL04o00r5//bOA1yKImvY66pIUHKOkiWJZBAkC0iQDIJkEQTJoGQBUVR0QQExfSISjAgG1pxWFwxrDuiaV1cE4woiKEj9962Zmtu3OdPT3dM9d67/nOd5H3Fuh1OnQ52uqnMO095dm9XWa5aw9fHHH6+jLU30JYJNVq9eraeZzP1Duph0KB8p2fPAVy9HNXeWxKORj0a3jMjvP7tLEyQ5uG4CjIBzWCVRLXOnUU+rYBNpf8mmuQFTjOS5lN6fzGDwt1RPQyZCsmcqYdp75MCuMZu5fXY7tWmcFuUjJZsmA3mgTy0bmb7OrT6De3Vyv/AzHUj29AO5Lb1W48ktKKYitcEPdh8wTziYQPofKp4Yo5x88slq/PjxavLkyWrKlClq6tSpavr06WrGjBlq1qxZGobwrcyZM0fNnTtXhL/Zt2edCMfhmBx72rRp+lycc+LEiTrXl9GHl9HIrk0DHYGSLmAyfPfeQ6rzWU20vkQCbt68Ofoop0527typ7UZ5yiDzb0lINk0FLOmgwoW5N0g4TEqJePLBBx+oli2zq2Qwmsla3twczZTs6XYE89B3H4r7W7HK0aNH1L6PnxS3s0LAjV2cAosMHJtzWEXazgptcCPpPIJJzsFW9arE7iveUUScgtXhZJt0yk8o2TNVMLVJRTNjG6/PLqOZrGnLzdFMyaZ+4eOjSTSfam73GZSnDDLPtIRkT7+Q/iffiSfE7o1081lwgBfNGBnovWr3AfOMgwlXj+uuChfKHzNQly5d1I8/JlgTFoKQHmDo0OwKQQzhzxka/Jom6QL6hZtoeP9IsBSdy/Lly6OtSb288847+kanBCVTCZK+QSDZNEyoWd+9xWlZ9jUP8F/VxRdfrPbt2xdteXw5fPiwviZ8rZv7qtlpldTG+UPEc4WNZE84cihR2p+jav/nz4v7xvgo5wgmcnDve/K2FqR0RfHSE1nh2HaJVzXIQBtoi5NgC2lfkGyaas7rGMnTCDiVpNgxwr/5zfydbaVj5AaSPcOG2s1jhnSPOd7JPrtd2zdT//7nRvFcYSPZ1A86+0U0h2+69BmUoMQPkPQNAsmeyUD/VqJY4dh9kS4+C0vV1l8/R9Q5Gew+YJ5yMOG2WQNVpdKRCjNAhQXWxaRKvvrqK9WsWbPY+UsULqhWTjpX1DVZpAvoF/JymZfnggULoq3JPeGrlOklqgVR71fSOVkkm4bFmql9c9yX5DFzGvmIJ/YRESpjLBndVTxnmEj2hF/+s0Md/SPnaKBVDn3/kbiflX2fPBndOluOHNonbmslXhS5tK0Vjm0XdJC2tUJb4gk2wBbSfiDZNJWwrMjM+JQpU0bMhcdvpUtHMhuw7U1pUi5SsmeY7HhojapdvVLsmQvq2S1VoqjactsS8ZxhItnUD+SfNh/L6dRn8E7cOC+cD2/JnsnyxpO35bi/cttnKV+mhHpuy0pR12Sx+4B5zsEE1oQ0q519wUqUKKGGDBnimWHDhnmGRKbmvKSdof6qpGMQSBfQD4xemvJT55xzjo6Atcr333+vy3qx5iWVcvvtt2udundsEcqUkmTTMKD+PKPYtAUnfvTo0ernn3+OttK7UIZtyZIlsUhKjjns7MYqlQmxJXsafvnPP9WRgz9FtbXKUcfUPQbJwUScHDY96nlUuD+zfnMajeSYkrhxMGmLNIpJ27GBtI9Bsmkq6dAoO2vB/fffH9X8WOFvZjv2kY6VaiR7hgV1mBnNMc9Z0M8u05DzpgxTP32QuilzyaZeYfTSlFlOxz6jRd3KoSwhkuwZBMQ+dGlnGZjKJZ+l2RmnqQ9e2CDqGAR2HzBPOpjAmqH+bRvEvrBSTacmNdW2peEmg5UuoB+oGU5tcfRet25d9FGNCB0MqTdOOOEEXdIrlcJLiwoPvNjvv3WxqHsySDYNmlHdmmr9sS1rbDZu3BhtXXxhmxUrVuipNSf5xz/+oSpUqBC75yg5maq1cpI97bD+0D7Kp6eNE0w/kxRdEqea4Dh08cTJ2YtXAz1hRZ6sNtiXA9BWt0FFkk39wjo4Ek+7vfZsmz9f5IOHcoZ258Aq/M2UPGSfRAmu6dS96uMVyZ5hsHjmKO0ApuLZpeQk72FJj6CRbOoVri21xdE9PfuMv6jFo7uIuieDZM+g4PpPHds/1l+kmqF9O6k9b28TdQsKuw+YZx1MQ5829WMG5MKFiTlP24bVQvl6siNdQD9YHcyHHnoo+qhGkq0WKVJE/z5u3Ljor6mVzz77TE971KpWMfCKGJJNg+SCHs2z7ovIPUFprrfffjvaqviCzc29RD3aRLJ7927VvHlzvT2wJiqd7j0p8CfRNHm8YCGmnfd9/IS4j7SO0ki89ZscK950fiJHUZoed+tcgmRTt9wxe7C6oHtz1bR2RVWySCFdN5x7hvVnBI+RaYASe9dO6KkT+Nv3NyX9gIX/iYRtzPbsaz3W/UtG6JyZPVrV0TM2RQrl19Pp6MOofdnip+jRpAt7tggsl6tkz6C5YvYFsecwVc8ua+DDmKmxI9nUK1YHM137jIqligZe8UeyZ9BcPKpP7J7gfgoTc57+Pdqm5N6z+4B53sGkhjMGZFE2X1PkKAsLvnI5FzVUJV2CRrqAfqCCTpHCkVyMJLI1wpA7vzVo0EDXRs0tIeINPYKsKACSTYOC/JZm9IOar19++WW0Nc7CtBL7wL333hv91Vm4Nh06ZNeRpjOXdAoSyZ7xOKayz9GjjqOK8RxM5OCed8V9fv85fk1e/ibtw7HiiZOzqEdLbaN+tFHaNh6STRNx59zzVIdGNXS0rLnWiSDHKs7mpvlDY8e5flLv2N+vvvrqaAviC9uY7W+Y3FsfY9XkPqpT4xqxpR9u4HloUaey3tfo4gfJnkFCfktSpaFzqp/dZXMvFHUKEsmmXmGUulCBSKW3dO4zgqycB5I9g2bJJaO17qn0WSaO7C3qEjR2H/BP5WC6ifhLRsgBxrnymoO5951tujY4uj/77LO6LS+99JK2WdWqVdUnnyQu4xdPjhw5op588smkXjbffPNNbBQzyGkkyaZBsGXJCD2yhD1LliypPv00ZxJvJ3nzzTf1frBhw4bor4mFdWH160dG6ynXRrCbpFtQSPaMx+ED30W1zJY/CNr56DFx+0iEtixHDv0s7pOzHnhO4W/SPhwrnsSNdM/SGd3tQhvF7eMg2dSJhSM6xzp0A/dWjx49dHoRUo9Qko/1cOXLl8+xHXBP9Durga4adcvMAbHfSWWSSNjGbM+0I2mL7EuPyAVZr149NXDgQJ3yhLyQjGBR+s9a4g9wNHu3rqe2+RxdkuwZFF+/sUWVL1tS65kbzy7leQn6kHQLCsmmXuHaURscndO5z2AUM8ilGpI9g8bqYKbKZ8k4mD7JOJiJ+e/r96uT8kVeFkTisY6lU6dOavDgwXoaJxm577779HHJ75WMjBkzRh9nw6q5Yhv8INk0CAi4QVdwCqBAfv31V/X888+r7du3qwceeEBdeeWVsX1xGLZs2aIeeeQR9cwzz+iF807CNF6+fBEnhEoskm5BIdkzHod++DiqYU6JV+PbaT0lYh/9jBcUZBV70I7Xcxji1UynjdL28ZBsGo8Zg9ppp8zcF23atNGjRvHW+fH8Mpq2dOlSnafR7AdE2FKu1oyCsl4tkbCN2d+aa5gptvbt26s777xTj4bEEwJbnnrqKdW7d+8c03JMqd+98HyxzU5I9gwKAm6Mfrn17PY95yxRt6CQbOoVlkawNAN9073PCLLsqWTPoMk4mAEhXcCgyTiYifnH1hu03oxCfPvtt+p///ufeuONN6KtSk6oZsGxmzZtGv3Fn6AP17BD60ZiG/xgt2cQbF06MpaLtW3btvrF6ySjRo3S27qBVBKJZMKECXpbHJLbLglvFFOyZzwOfP1aVDu7HFW/fLnzmO0TOX/2SkAH/vtq9C/xhW2s+ySqxCM5mOiKzpLQRvv2Tkg2laC+s3HqeD5XrlzpKTKX0SA67Dp16uS4l8wIJKOdTsfjb9KIKPn6Xnst3nWNL+TXtDq9VcsV16OqUtvjIdkzCPa8tTWWkzA3n12m598McRRTsqlXWCoR0TX9+4xGNSuIbfCDZM+gyTiYcWjWuKEaOXyomj93tlowb44aNmSwuJ1BuoBBk3EwEzPtwsiUGS/BRC9Vr7Jq1Sp9bNbkJCPo1a5du6zO9nj17rPrxHZ4RbJpsiwY3lm3FxKNgCCsbzvppJP0i5p71DrCw7/5jb+R1mTkyJHRveLL+++/HzvG8C5NRB2DQLJnPPZ9+kxUu2OF6Wt7ve94qYOMHP3jsNr3cfY+TvkojVgDi9iXYziJPSUSOjpNw9NG6/aJkGxqh8T8ZYpF1khxTRkp9CuMIl577bU5kn0bnAJYrNO+ULx4lkPocn1hPCGR9FlnnRU7JpVgpGCkeEj2DIJNaxbEdMrtZ3fB1OGijkEg2dQrA9qdrvXMC30Go/XrZgdTXleyZ9BkHEwbjRvWV507tFOLFsxXN6+9McbUyReL2xukCxg0GQfTGdYclSweifq74YYboi0JTsy0ESMCycptt92mj7Vw2gixLV6RbJospMZCRzoVvurdCFOdv/zyi+54n376ab0/8KL94Ycf9FokHAQ3wkuVNVDsTy5YSccgkOzpxNHD2XWa7fLbT5/n2PbAV69E/xJfDu55J7b94V/2Rn+NL2xjtmffRIIOZntAx3hC26zbukGyqR0+EMy9QNWYIOS9995TdevWjR0XFi1aFP1rTuH+NSmKoFGjRmJCdj/Cu7hJk+z2eQlMk+wZBKSIQZd0eHbJiSjpGASSTb3AGnOyBaBnXukzRgT0sS3ZM2gyDqaNIYMHqhtW/E07lTfduCbjYOYhB5MvZXRmZMLtS9WLmPVbLPxPVvbu3atHDOrVrhpISgXJpsliElhTZs+PvP7663p/WL9+ffRXb0KgB/sz/SjpGASSPZ04vH9PVDtJjmY5dC/HtnXjYB45mF2G8eiR36K/xhe2MduzbyKxOpjoho7xhLaZbd0i2dQKo5cmDQwl8IJ8Ngkq6datW+w+Ywqc9DJWwXFiGtxsQ2efTIJxSXBWixaNVLeirSwvkWxhR7JnEAzqFYnmTodnt/5pVUUdg0CyqRfMh09e6jN4FwaRvk2yZ9BkHEwb8+fM1g7lsqWXq4vGjVVr16zOOJiCLkEjXUAv7Hp+fSx6nOoSQcvXX38dm5J7+OGHo78mJ0Slsr4wiDVKkk2TpXX9SP1mokL9CDV12R82bdoU/dWbDBgQWfJAaUpJxyCQ7OnEoe8+jGonyx+/H4jluHSzphL55YsXHVMa2YVt2ceNmDWb6IRuTkLbrG11g2RTKwT2mPuAYJ2g5bffflP9+2fnw2Sk0hq1e9lll8X+1rhx49DenZdffnnsPFS8kmxhR7JnEJzbtbXWIx2eXUoHSjoGgWRTt6yfe14sejwv9RksPQhiTbpkz6BZMivjYObg0pkz1JRJE1WbVs1Vj3O6qBtXr8o4mIIuQSNdQC8MPjfyxV62bNnARycIDjjvvPP08VnU73aaKJFcd911+phXzx8ntskLkk2TxYxgYlM/a5OINuWLmxciaT/8iMmrl04jmG5GJX/735d62193vxH9xVl+++k/6tdv3oz+X2JhW/ZxI+iALuiUSOzT6W6w29NOmwaRqVLeW/bRxaAEJ9M6SkkOQ+5ZgneowsJvjJ66zQPpR8jzZ9YdUv1MsoUdyZ5BYEYw0+HZTdcRTPKwGhvltT5jXK+WYpu8INkzaDIOpg0cyyZnNND/zjiYecPBfOLua7NsEnmx20t9JStMr7FmjGPzsvWSEy6RmFGCti0biu3ygmTTZCGptbnfvvpKLkOYSGjjjh3OgS7xBNtTxxYdzqx/qqhjEEj2dGLfx4lTCSGMHLp1MAnU+d2FA2iEbRMF9xhBB7cjqbRNarMTdnvaKVciEs1M9HeYwhTnaaedps8FTO22atUq9v/btm2LbhmemJKJNSuWFG1hR7JnEFw6MZIkPB2e3V5dzhR1DALJpm6gMpT5GMiLfUbD6uXFdnlBsmfQZBxMBzIOZvo7mD/uekQ1Ob2W1rVly5Y6lUlQwhQH+dA4Npx//vm+RgPiCbpWqlRJFShwkg5QktrnFsmmycJL2LQ9jAXwiYR8g+b8k/q2FnUMAsmeiXCKwjbyx+GD6uDe+BV2jhEv95aHbdEBXRJJvCTuiZBsath+1ZjYNCRr8sIWOuD8+SNBGyYXI5C3MhVC8BDnK5/lVEv2sCPZMwj46DZtz+1n9/olk0Qdg0CyaSKI8q9VqZTWLa/2GVSdIkBJap9bJHsGTcbBdCDjYKa/g7lm2VStJyk0Xn6ZAIbkhRcC6UuYOuHYQGUPkhEHLUOHDtXHf3DdFWL73CLZNFlwDqgegX5EhB48mNhJCUq4Bqw34twF8p2o7rnMW35BL0j2TMTv+76Oauosx5SWzAVxqwNtktqaCMmmBquDSTBOKuSqq67S5zPwviTiPBVSrVo1fU63SzokewbBTx9s19XCtC65+OwWKlhAffHqPaKOQSDZNBFTB0TSSuX1PuOKC7qJ7XOLZM+gyTiYDmQczPR2ML956wFVrnRxrecFF1wQ1Tw5IRq0X79+sekTQ4sWLaJbBCs33XSTPv6M8YPENrpFsmkQzLQEaFDCL1Vyxx13xM5LnjpJt6CQ7JmIg9/uimr65xHaJLU1EZJNrVQoGUkdVqNGjeiZwhXWY9auXTt2//Tq1Sv6l3CFdYs4LZyTdaeSLexI9gyKW5bPjNkgt57daWMHiLoFhWRTJ8hoULxwQa1bXu8zBnVoKLbRLZI9gybjYDqQcTDT28FcvuAirWOhQoWSDh44cOCAjgI1BfOhYb3qavR50VQbPqMxEwkjKxy/RaM6YhvdItk0CBiBalCtnNaRFygvN0mYuvnwww91SblrrrlGTZ06VQ0bNkxHkhLhy1QR65KuuOIKddddd6m33npLHTp0KLp3TiEHn4m+LFP8FF3KTdItKCR7JiJSCefPJVIlIjdINrVigsW4f5Kp6+xFbrnlFn1OSCapuxe59dZbY+ec0LuVaAs7kj2DglHMNs0juWxz49mtUrGMLt0r6RYUkk2duOjcyJrcsPqM6hVKqHNaRNYBh91n1KlSRmyjWyR7Bk3GwXQg42Cmr4P53XsPqcoVymgdL7nkkqjW3oVoP2rvmqktKFbkFHXN/PH6HCsWT9S/nX766dE9ghUWhJcsWVIVLJBf7Xl7m9hWN0g2DYoN84aoUkUKaTvQUc2cOVNP/Xz00Ud6fVfPnj1VsWLFYvZzCy95qlOQIuRf//qX7ujoBM0auvz5TlArJ50r6hQkkj0TQTUcFeDaqlyXrLbYqxC5RbKpFeonm2ueqpE0UwMa+HfYQpSwGTWlHObmBUNFW9iR7BkkH7ywQVUoF1lvmMpnl/fZc1tWijoFiWTTeDx05ehYNamg+wxyn47v1VKfY2KfM/VvYfcZvB+3LR0lttUNkj2DJuNgOpBxMNPXwXzojkiFBFJp+I2SZDTFmtqEurnD+3dRH+3YFDvP5ZeM0X9r3rx5dK/gxaxXevrev+VooxckmwbJrbMGqLLFI/cE8NVOh2X+38AUIelgiBim9Frr1q01TBexJolE2FQXse8HvDTNvwsVyKeuurC7qEvQSPZ0w5FDwaY2yU2hLVIb3SDZ1AqdbsnoB0rBggXVp59+Gj1reJJqB5NSi+Z83ZqfJtpBQrJn0Lz+xK3q1ErZawPDfnaLFC6ktm+4StQlaCSbxuPKsZHZqCD7DLKXdGlaS22an/1BMaZ7c/23VPQZf5vYK0cbvSDZM2gyDqYDGQczfR1MM3XN+ioWWK9evVqX0uLfboRpM1N5A5o2rK2euudYB4+1kfy9e/fu0T2Dlzlz5uhzXDXPfz5MyaZBQ6BNq3pVYjYDbEiE7sqVK9XOnTt1qhina8DfKEdHXWimMZl+o+OyHrNWxVKBJBJ2i2RPN3hJK5TuQlukNrpBsqkdE1gB1O4OKi9gPEmlg0kqHxOxfnKBk3I4G4mQ7BkGn79yj+p1dnbKJgjj2W3coFYghSPcItk0HmbqOqg+o3alUqKDx9pI/p6KPmNcz5bHnN8tkj2DJuNgOtChXRs1fepkNWv6NDVk0ABxG4N0AYMm42Bmw/pI9OMlsXnzZv1vvspfeOGFaAtk4WXCuhnzBV+qRFG1+sqp6oddD4vn6dOtjd5uwoQJ0SMEL6x94hwkR5Z0cINk0zBYO72f1hVYJB9EdCrTa9YRoDlDO4rnDgvJnm44uMdDCqI0F9oitdENkk3tsJb3jBrZzgj3jtuO3Y+kysH897//rUqXLh07l9sKPgbJnmHx8va1MT3DenbXXz9HPHdYSDaNB+sj0THZPqPoyQXU1P5nqYeXjRbPYwoLpKLPYH2zpIMbJHsGTcbBDAjpAgZNxsHMhjU+6PfII4/odUT8m6mPd9917vTXrs1+ybIA/sMXN4rHB2qE16waSfXBAv6w5OOPP9Yvrzo1q4h6uEGyaRhM7B1ZX4S+H3zwQbQFyQvrwsxi+R6t6ojnDgvJnm5wm7xckt27d6vnn39e3X777WrhwoW6w2fEg+lI1vJVrFhRr41jrRvwb37jb0y9sS37sC/H4Fgc06+YcpJ+kGwqsXH+kNhUOUycOFE7KGFIKhxMgi1MYnXo06a+2G4nJHuGxd8WRdaTh/nsjh3aQzx3WEg2jQdrFtExmT6DgMeN84aIxwdqhFcsFcmakIo+o0qZYqIebpDsGTQZBzMgpAsYNFYHkzUkP/74Yyj89NNPsRdGujqYJ+WLrAX6+9//rurWratvrkSVOljYbhahd2zTOGFQzdtP355l6+P0g8xIRVjCdGGRIkVU/pPy+Y66lGwaBmaKvHLlyo4jUPyNxfA4EMC/E41YkYibY5PWhhe1dP4wkOzphn2fPJnV0D+i2seXPXv2qK1bt+rAgo4dO8YqnIQBx+YcnItzcu6EktUG2iK10Q2STeOxZmpfHRBh9O3bt6/njod76bPPPlOPP/64DixZsGCBGjt2rD4WSa7PPPNMnRLJnINo3nPPPVeNHDlSXXrppTq45cEHH1S7du3SKY38CInErcExlB1klFZqsxOSPcPCTJGH+ezWOLWC/jCXzh8Gkk3jceIJkRRSfvuMxjUrJAyquf3SQbq/SFWfkS+rTX6zbEj2DBqrg5kqnyXjYPpk2NmNtQHB3MRhYc7To2VqRpOkC+hE1cqR1Dk333yz7lTefvvt6KMXX6hPzD4Vy5dylfzXBPgwasRLNkxh5IpzPXu/v8hLyaZBQ7CGcQ5Gjx4d1TySd5B6xcuXL1eDBw/W0ZMkHOaBJ2UJMApHAAEvdtZALVq0SD3xxBNq//790aMovT/HPu64v6g7Zg8WdQgDyZ5u+e3Hz6LaZwspXHB+SPdCcAQvV9oVD0ZRSIaNY4Rthg8frsaNG6cjfq3wG39jG7ZlH/aVjmngWUYHdHnsscfE9DK0QWqbWySbOrF6Sh9V7JRIKhugvCORyPEEB3T79u3aaWb9ZuHCkdKTQYDz0LhxY3XRRRfpFDyJHHIcrqVLl8bqm0OXZrXiTpcmQrJnGHz//kM6Owb6hvvsHqfee+4OUYcwkGwaD1Oy1E+fUaroya6KPZgAn1T2GSsv9pdpQ7Jn0MybMkzrCFb/IgzMeS4YkppRdLsPmKcdTL78C+XPLn2WKvhCWj6+h6hTkEgX0IkRAyKRfG3atNELz+1CyTg6Y0Y6kNdffz2WBHnDqrniMa2wJrNalciaMV6oYQvTnZxr7VXTRX0SIdk0aFjQjo7A4vj7779fDRw40FeaEwMdGBVemOZlZMH8PqV/G1GHMJDs6ZqPHlOHD3ynryG5BAcNGhT7kraDM0OngDNz4403queee05/1ScaHXISOjGOwbE4JsfmHGbUxQ66oSO6IuhOG8S2uUSyaSLWZX1AVCufPZKLw4YDaUYzCTjhnujatWtCJxpwglhCgDPdtGlT7YATAc1yApymU089VTum1o5Igo8B9iEf5Jdf5gziev/99/Vxs7c9To3o0iSp0XbJnmFAhgqjd9jP7qorpog6hIFk03jwIYB+fvoMUm1Jx7TCRwYlQtk+lX3G9IFtRX0SIdkzSHY8tEYVPiV7SUyqYCbwsc3LRZ2CxO4D5lkHc/2cwbG1S7wgSX47YsSIUDnvvPNiDxejVrfMHCDqFhTSBXSCFyYvePQjAbC1k6aiRs2aNfXfrr32Wv03M4VzRr0aOgGxdEwrt103S29P5/b5559HjxyeoCfn81v5QrJp0AzP6kzREawjOIbixYvrFB6TJk3SozxMRTJaAKtWrVJXXnmlmjFjhp6uxBmw728d6Wt7ejVRhzCQ7OkJnMxf9uopWmt7TAfM6A4l6eIlpw5DOBfnxFFCB3Sx6oau6JyscwmSTd2wdelIPUPCiLXRi9EzRo0kJ513H7kHcZC5l1gCQNJvpscYWUwkOOOMurH+EIeI6GlG83BAzbvOCvc49yqj0bNnz87h6BLosXRMV7FdXpDsGQYLpg7P0S7zb0OQz26/7m1FHcJAsmk8+EA2Hxhe+owaFUq6Wv4wa3B7vX2q+wy/lc4kewbF+8+tV+XLRlJX5YbPUrzoKeq1x28RdQsKuw+YJx3M+xYNV6eWzf7KZFF/quT666+PnZcvs80ukwf7QbqAiTi/XyQXGDcwnc4rr7yiR0D4N7+zHu2bb77R1SXMi+XemxeJx7LCOkiqULA9FS1SIawJ43zndGwh6pQIyaZBY40CBmzKaBEd0muvvaYTALsVOntG0ei8mK6yd3olChf0tabND5I9PZPlqG29Z512VsaMGaMefvjhUOoQ+xV0QSd0Q8cH7r49EOcSJJt6gfyEppykHRxNRtrWr1+f9Givk7COi2dw/PjxOepJSxAlHNS7ULJnGLQ/84wcbQjz2S1fpoSrj/ggkGzqROcmESfSS5+xaOTZ4rGssA6SqmNsn+o+o0WdyqJOiZDsGQRf/us+Va/WqVo3yC2fhRnIT3ZuFnUMArsPmOccTNa8WTt1FqmH9YKNJ6zdMuenNFUylQOckC5gIva8tfWYFyeJnM2Lga9v1hjxIuX/iRpP9OJjgTrJ1s2xUlXajuk39GaRvKRXIiSbBk3VcpG67wbWBDKVmayQLoVRPusoEgvyuf8lPYJGsqcf9n36tDr6h/uOOrcEHfd98rTYBj9INvXKg1eMUkUKZU/rt2zZUm3YsCHHOr9UCc4W61X79OmT454sX7KwWjyqi6i/XyR7hkG92pHUOYYwn10CMFnzKekRNJJNnWDU3P6h7NRnEDWe6EOXJRIkWzfHSnWfwceZpFciJHsmC9Xv2rXK7pNz22ehBHMyFfKcsPuAecrBtN60cPbZZ/uOeExGmHpiWsTo0a5h9VBGlqQL6AZuaBYSFy2cc0rtjDPO0OtsGLHh/6nS4yaA5tqFF8VeNkyjpEqoa8vUysmFCqhv331Q1M0JyaZBs/yinnq6yGpnXqgs/F+zZo1ew+QmgTYjIKTZuOOOO9TQoUOPWQfGSMDsoR1EHcJAsqdfft3zjm7jF198ode5kSLHDr8HiXQOCXRC0FHS3S+STf1glgGxBtKpU8IBpBNnmpv7bu7cuXqqm/dUhw4d9BpUAncaNWqkK9K0bdtW9ejRQ48sESy1YsUKXeqP9DSJckFOnjw5dl+GEXgm2TMMHr9ruV4eZNoCYTy7zPzcsXK2qEMYSDZNBB+uBMySFN+qu73PYAmWmwAa6pubZR650WcUOOlE/YEm6eaEZM9ksA7OQLr4LAN6tgtlRN3uA+YpB3NE18gXFLA4nQhHXqi5wT333BPLMQUsbJd0TgbpAnqBae37blkcG9FkzVmZMpFpbpg6tr+4n5XNNy5QJ0ane7hB3azrCkp4cVepUkU7t7ueXy/q54Rk0zDgw2fZhefodEXUXDb2NTClydc/05qMklx88cXqwgsv1OvqyN1Ipy8FFtDu+lXLascyVSOXBsmeyfDrj1/lKJ2XLqDTgR/8V+yJh2RTPxgHs1WrVtGnIiKMtDG9j3NIkI31XZQsdNANGzbU9+rGjRvV119/HT1rRKZPnx7b9s6554l6J4Nkz7DAAXjkzmWqZ+dWKt+Jx67D9Pvs4oi1blZfO5apGrk0SDZ1C9PajEibEU17n9G/bQNxPysLhneOvQdzr8/4i1rv496U7JkMl00fEbNduvksC6eNEHVOBrsPmGccTAJqTABLOoJu10/qLeruF+kC+oHE6eVKZ0/lMnKJc/njrkfE7Q2Pbrom6wUT+aLlRRrE9JFXIeqV86OLpKMTkk3DhnVoE/ucqfPDnSR0WIngxXxa5dJqVLemKS0NaUeyZzL8+u2HqkGDBmKbcxN0QjdJ52SQbOoHq4PJmkjKETIKYg2ukeDjhM6Ezpb1pYxgks4IOBYjU9WrV9dl/qRgHisEqzRp0kQtW7ZMj/j+mRxMKx/v2KxWLJ6oyAds3nte4EO8eaPT1OKZo1JaGtKOZFOvkDi9eOGCsbbRv+FcPrLMeabumvE9Yu+93O4z0EXS0QnJnn4hoIa+1tgw3UC35x+4XtTdL3YfMM84mCwqloyUTkwbcJaou1+kC+iXT1+6Sy2aMVJNHtNPPbcl8bQ46RTMFDu5Be2jGKkSavuiw7oV3qeYJJumEtY2XT2uu6puST1DZ03UL9GZplYz4EjMH9ZJB7BJx0o1kj2T4fD+PXpq6NNPP/UE6VHcIu2fCHRCN0nnZJBs6gfjYOIsknbI3C8GHEkSqBMtSnlCghyY5qZjZzQnkTDtzhQoybOJDCdIhVQvOKBSZDXOqHUk+s/kYFphLfvfN16tTq8bKb8L8Z5dIoM3rZ6vAzmkY6UayaZ+uGvh+Wpk16aq31kN1MpJiafFSRtoptjToc+YPcT7kiLJnn4heNbcI+nKjcumibr7xe4D5hkHk87XGIX1ReS3SwdIeWL0urhva1F3v0gXMBW888w6HfVIm6gpHGQJNa8yZ84crccVs73bQ7KpX/hyJ6kwI+m8SEmMfeO0furmGf3VrbMG6NFG/ktdcr6cSc9BxacyxbLXweIksO7PCClzrGX1ChfKr7o2q62mZn2oMOXOeTifOTbn4vj8Dvz/pvlDfSe0dkKyp1/2ffKUOnokdemIvAq6JVO1R0KyqR+Mg2mF+wiHUpq+DlJwUikhSP3o8uVzBoEY8oKDyUzN56/co0eUdj68Rv3zwdVq5yM3qlcfvVm9/sSterSR/760fa2eKSEdG5VPKlfInhpO9OyWKFZYjRzYVa1ZNlVPuXMezmeOzbk4Ph/uwP9/tGOTzi0s6ZwMkk3DZt2lg3SWC2yRLn3GBT2ai7o6IdnTL3x0mPsjXX2WlYsvFnX3i90HzDMO5jyLg/nmm29Gb6Xcl71798b0YmGzpLtfpAsYNqzbrFszUvqQlyov0twUk2LBzXpRO5JN3YJDed2Enmpo50Z6PRJ5T625Cb1C3kUCAezy3Xff6QX0iaYp44FOLGivXamUHmkgD+E2H4vb7Uj29APO5W8H/qejO72kfUmVoBP1sw/u/17t+/hxsQ1+kGzqB+s0JWstN23aJCbEDluw05NPPqlz91lHNtMxyAeH8sl7rlNzJg3V0bvk/zNBin4I79k9TgcwNm1YW88sbb19qdr7TvLRvZJNw4R1m9T/pk3p1Ge4WS9qR7KnXzaumhe71unqsxDAK+nuF7sPmHEwk5Q/k4PJgvf+Pdrqtpx44onq0UcfjbYy94RF0egzqFcHUWcnJJsmYuP8IWpIp0a6DJq5rn6g06lTp45er0ZeOauQf/Hnn3+O/l9EqNG7ePFiHS2M7aVjugVnuGerukkVApDs6QcSlxNZi15MrRK1jJOUW9NnCOdm9A9dzHQvQRuHvgtuLaZkUz+YEUzuCych2pl7iBFHEoJTAYhEy0SKEzFOoAqBO6zHZD0l69RwnGj3tGnTdFodou9J0k4krpNMmTIldq+l0wjmv/+5Uc2+eIgue2v080NuPruUrrzw/J5JJcSWbBoWBDi2bVhN655ufUaHRtVFnZ2Q7OmXjIOZBxxMRpKYApwztGPMKNTo5YWaDtBZGb3G9WqpdU2mTJoV6QKGiXVIn4oe6SDPPvus1qdbh+aizk5INo3HfYuH6y9ee2AOFToolcbaNNK4UG+YEoQvvPCCevHFF9WOHTvUzp079Vc7UEqNEbEffvgh2oJs4X4hpxxTSKRDueyyy47prBCSHO/atUu98cYbuoPjuJyDc3FOzo0OjCix5o7AD5JhU+vXOlJz/F//qjo2rpFr0ZS//GeHbg+5E602BfRkLRs54UgJQ9tMScQghWNybM7BuTinNJrVu3dv9cehfWI7/CDZ1A/WIB+rEPCzbds27RySH1Nan+kXHIX69evrtZh33nnnMeUh0y3I56vX7tMzHPbAnLz87J6Q5eSe17tjWmfPAOvStXTrM5r7SLYu2dMrjKCz9GH99ZGpekhXn+Xq+eO0rgwuSW3xit0HTGsHE4eN0Zj8+U7QSaaNUagpzEOeDljLzdGhM11Z7JQCOqeY1CYvSBcwLHgoalWLlDvr2bOnqwCBVMjbb7+tdWrZuK6otxOSTSVIy2HWDwHXdOzYsbpjSNYO7E8+PUY4iOg15zBQjo4Om3Px8CcrTEVfeumluvqGOUfBrHtyUt/Wnj58JHt65bcfP9U6Mepz991369Eyp1RFdLA4BeRtJIcjnfhNN92k7r33Xu0c0EEzEkAQC/BvfuNvbLN27VpdIYN9OQbHkpxJA7qgEyMe5H48euR3sR1+kGzqB6uDieODPTp27JgjyESCgBTSohCUQjQv0+vt27fXUHeaUUycbe4/KZjHCsci6IcKNwRTpZODSRo2s14c/mzP7iknF1TXL5nkyQGQbBoGDP5ULFVU65mOfUbdKmVEvZ2Q7OkFHDZGoQsWyK+T65vrmK4+Cx8yLNMoU7KYmj91mNgmL9h9wLR2MOtVdS5Pls5Ur1BCbJMXpAsYFkRMojejF7m5QNsulMLDSahdvZKotxOSTa3gcA3ueEbMCWFqjBx3//3vf6NnP1aIumX0CAeH0mlbtmzRJfsYJSGKd968eToRNdOTlIxjxMN6X7Bm8vTq5XRpPXvarSJFiuipS6aUybfHYnVSw7CmaN26dTrIAGeK0ZFvv/3W8YXO6ArOlvVlQi1zt1WnJHt6IRLYc2xCYXSmDN91112nRzYTlSAMEs7FOTk3Ohxjv6xru/+LF8T2eEWyqR+Mg0k+RjoHe5tw/mrVqqUjZ6nDTG5MRtAYSXNbLYQPACLqn3rqKT3SS75HkrJL0708I1YHKLccTByuWRMGx56h1Dy7x6mzWpyu+nRrk3W+nOlnwn52+3Vv67r6imTTMCBDBrqla59RqXRRUW8nJHt64cymWU5V9JrlNRrWqy62yQt2HzCtHUzyAdLwUqVKqc6dO+cJTGQhX3ZSm7wgXcCwmHJBP603efLSSXjZ0okS0Snp7YRkUytEe5uHiylGRiIkoQ4vHS9Jg4mmRR+zn1sY2e7QqIZaYamCQWR4rzPrqqInZ3ckbuEFyggc9xwdmRSEgPC7dfRlQm9364Qle3rh0A8RfRKt50PoELZv366jGwmaaNeunU5zkijXowT7sC/H4Fgck2NzDifB+UBX1oxK7fGKZFM/SFHkODM4Moy8cm+GJTipJGieNGmSHg226wG55WAS7W10CPvZZYRn8Lkd1DP3rYidn8jw8cN7qVIlIiN4XvD77F532YQcNoiHZNMw6Nc2ktc2XfsMMnhIejsh2dML5EHFJnnRZ2EGU2qTF+w+YFo7mLUqRRZr83LIK8LXPzr7rYVqRbqAYWG+vFJZ1suNMHVJB8I0mNfSVpJNrTCax2gi7QaqdRw6lJ1O56WXXtK/OU1HMiLJKEqBfCfqutGls15qjF6TaL1Ls1pqTPfm6qoLuzuOHLJul/JrBIn1aFlHNTutkqpVsZQuD4nziXPK8gunKHZeqEydEuRhRkdwmhYsWBDbhhfuOpdRv5I9vfD7vt3aAWL6lTyNpOl49dVXHUdu7MK2TAt/+OGHel/WrRFEwGgQ8G9+429sw7Zej8++jDahI7pu3rRRbI9XJJv6gVrf1utMYvjcGC36/vvvj1lLy31PYQFJ72SQ7GmH0TxGE40u/p7d4/RIZKGCBVTJ4kVUpfKl9SgOidZHDOiiLr9kjNq+4SrHkUPWr1Fud/mCi9QFQ3qoru2bqcYNaunykKVLFtXOKdOQnEvSAdw8u3xgv/vsOlEHO5JNw8DMMKZrn8GyJ68lnCV7eqHJ6ZFS1nnRZ6lxagWxTV6w+4Bp7WDWrBhZr5VxMMOF9Zem0g9r2dJJKDPG1CYva68l1ySb2tly+QjVsHp2jr8uXbroNTwEfVg7hXwnHK8a16qo19bOPb+jHon8v0sG6tyYOI+UcgwquMsODiiph0jCTlqYGyb3VgtHdFajz2mmWtc/VRXKn7MTpWoLwQUTJ06M/VaxVBG1fo77lDKSPb1w6PuP9ZSjVS/gWjIFSfAI6/lSLZyTc6ODND0/d/YssT1ekWzqh2sn9FRVy2VX4QIcYSLAaQeOX1jC1DlOD4EyTNFbdWCd+YxB7USdk0Wyp8TuN7eoti0bxnSK9+zmPymf6pTlNM6bMkzdecNcPRL51lP/p7549R7tPPJeCSrIwQ4OKKmHSML+3nN3qH9svUHdtXahWnLJaHVu19aq8Ck5R6ilZ7dm1Yrq/efcB/tINg0a1l8Wj65bT9c+g49zryV2JXt6oVH9mtomGQczQp5wMEmvQQRfXoDpAnSmQ5fa5AXpAoYBL1jzonvmmWeit116iHlZkMj4u/eCdzABB7FF3cq6/XZKFSmkLuzZQjuS0r7pAPrT2VsdEWsHW618CZ2QXdo3HpI9vcAazAP7f9KBNzwTrJEz+lgpV66cfhkTSLF161Yd6GAdifIrHINjcUyOzTk4l6QDuqEjuv68e5fYHq9INvULHxhcX9aU2XXH2SSKnOAQIqU/+eQTX/lGGTnbvXu3ruZDMA/OmhSZTqc9omtTtWXJCFHXIJDsGQ8cxO4dWxyjJ1QoV0otm3uhdiSlfdMB9L/5mhmqXu2qMb2tz26DOtV0QnZp33hINg0aHDfzYZuufQaFK3LLwcyLPgsfMlKbvGD3AdPawaxTpUzsQctrkHhWapMXpAsYBnxlk4wYvZmC44YLCnLwsR4OiGAlupfpIGAhPWtAqK0MjMow+sDUFmvMWLRPlC96MYUVxgimgRcRVXTM9ct34vFqRJcmjlPb6QajCtMHttUvVtMOksSTgkna3gnJnl7Z/9lz6sjBSC3iPXv26ICKQYMGOUaSAw4fa/6InO7bt6+OCp41a5aOKmdNJTkbgX/zG39jG7ZlH/aN59Aa0AFd0AndkMMHvlc/f/SY2BavSDZNFqb7SKR/1ulVHevc4xjWrVtXP0+kZiKVEdOtOI5MZ2KzmTNn6jREvXr10gE9xYpFEmVLMBXOUhKc3FQ8D5I9neC9QBUdo2+BLMdn4bQRjlPb6QazSGuvmq4/pE07SBJPCiZpeyckmwYNHz1keEHPdO0zWLKUagezRaM6seuX16DAitQmL9h9wLR2MAmAkAyRF2jhIweXHekChkWb5pEF2+lK2VLFtSMs6R4PyaZOMMU9rmdLPZpJSUZpm7wAo5WdmtTUpSq9vmANkj398aj65cuX1G8/fa7++P1X7cgxWkZCb8qWMf2KM5QoVU4ycGzOwbk4J+c2a93QCd3QEV3lNnhHsmmQMILIUo2zm9bSa3WTqTIlQed8Zv1T1eR+bXTxAUmHsJDsmQimuK+aN06PZr68fa24TV6A0cqhfTvpUpVeZ2wMkk3DoEE1eUYgXSh+SkHtCEu6x0OypxfGDesl6pIXOCfr2ZHa5AW7D5jWDiadI/WWKbTPWiSifkmNQJ3mK8dmc8UF3Txj3d8Ox+c88UCPeKAnBDGlKl3AsGBt0EUjztWL23nBETU5sFf7YxjQs50jVAKyYv+7/XhU6LHCeYEkwzCkTyfN3xZNFPV2QrJpBndI9gyC/Z8/rw7ufU8HAR09nD0VTgQ3KVzIl8koGyMR3bt316NrlStX1pHTpEOxTh/yb37jb2zDtuzDvhyDY3FMayQ75+Tc6IAuko5BINk0THACF4/uokZ1a6o6Z31cNKhWVpUrUVjnQLUHiJnANEZBWQJCtg6qsVAWFaeV2vdhrSd2g2TPDO6RbBoGrAU/t3U9HczIBy1ZMtqfUf0Y2jV0hnvPiv3v9uNRoScnNTQUlYBOUSb2PlPU2wnJnl5gNJ06889tWameuPtane2AFIDUp394/ZUxHlx3hWes+9vh+JwnHugRD/QE6vVLbfKC3QdMawfz/3ekC5jBPZJNM7hDsmcY7P/sWfXr16/roKDD+7/R1XSOHj0SdQdzCpG1BJ5Qixv4N79JwjE4Fsfk2JyDc0k6hIFk09ziwWiA2N0Lz9fcuygSmCZtmw5I9szgHsmmGdwh2TODe+w+YMbBTGOkC5jBPZJNM7hDsmcqIUjoly9eVAf++6r69Zs39YjjwW8/0M4iOTY1Wf/mN/7GNmzLPuwrHTOVSDbN4A7JnhncI9k0gzske2Zwj90HzDiYaYx0ATO4R7JpBndI9szgHsmmGdwh2TODeySbZnCHZM8M7rH7gBkHM42RLmAG90g2zeAOyZ4Z3CPZNIM7JHtmcI9k0wzukOyZwT12HzDjYKYx0gXM4B7JphncIdkzg3skm2Zwh2TPDO6RbJrBHZI9M7jH7gNmHMw0RrqAGdwj2TSDOyR7ZnCPZNMM7pDsmcE9kk0zuEOyZwb35PQB66n/B6RKNpFsW4FvAAAAAElFTkSuQmCC